��/  ���A��B�c�qG[��I��0*p���#漭l��������h��/�n����$�1�a�~��/$����}uXzyh����>�k�X��C�̠�����x��A� (=}H7Wc���4j�T�	�g��/1�����,�<k��B�bѕOev�$��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�UtK��^�)A���Q���=�.m[�F|��]C�9o���m����T��i���`3��.uFh!%�S)|cph$��ڞكRy�4��Ӌ%����?;� ɞ��8������ ���$I�.���_jbsG%$wm�G����J�A�&�ɇ�!�1R,Yy��fQ���h��*��Ӫj��H���G�*��<5 H�J��E��g�]B�#Gm�������P�Pglˣ�v+�ȇ�M���JD�'x�9KY2˒-�K^�B_�7�HE��	$�usfƩ8��0c����mv��g�t
�=[�Fg��:ql�ܽ�E�pz%	~,�-{d��M5�D�b��]�$~��J�M��f�}
�Q����Xhn�hw��ɻ�bw�}Ӣ��{�!x�UB\�]0���RDK�|1����0�E����!Ej��Xy?:mWu$҇<�;�_��k�$�R�N3���F���du��A���UoW�X/ #�J޼��L��t@q�5����UϪ�c�9쫃�#��{|P��+��q"��:A�#>�:~�">!z�����v�
"k<��J��zi��Gs}�U�Դ�����_�$-9����1�(�jXO���@)����x򮥅�-o�sm��ӄg�*��,`m��2wA�ގ�O30m�p��µҮ�4�ݦv���L$��*��dئDA�Rl�����j�T�C�P]�b!����P�kU��[Q����c���罆�P���UH���?��f���*�;I���Z��������6(Yǆd�r,+�&����=>Aţ�K2!�1�u̮���ؑ8hi��,�:����Mӟ�y9A����6�.5�u'Am��B��op�������e�N��{����Q28Bǻ���Jɇͥ;, �W��'շ �'��<�$9�-��J�ªQ��u ��[�kpl�ݘ��*N<ih�nE��Mx_�ɿ=Ć�"5���No�3ᜓ�Ō�a�����Lr�D�]�C�Z��^r5Ifs��ؾ�+N��B����~+�vC��ͺ>!d��d��vsǝ C�0����YD����n����!	����@��W{{wv��A�kױ�Ƀ���%%�"�LZŤ�'�Q�R���1��K���qxEG;�>S�����[0��õ�b�cw!�_ץױ����R�����(# �
��xa�����$���]
�A�;�)��z���<ݛ��צW~u&��`R�k�s~p��pT����6���=�g�-��Ə��}x@E/��5�P�w�^�Kv��FMR�y XL�7?&�fS� #ȕx]�D}Ň�pX,ࠦ5@��GHhf��&&Iґi��OJrK�r�4ޔ�Y��1����I� �ݭ�0���ߘ*pO ��3��0��j�aqG��R��Fh;)7W�P/����)M��\�y�����_��>�ƨA^3��YU]3I:��v@���^����3��>�4��#�R8� MJ%AK��''�N}-(��͊�֚۝fn���v��V����}g�����3o��9I��]������R:�5�=���BM=��C��P�ڵ�sХ�Ι�\1n\�7�f���
�Q�%V���9��sI�qQ��L��Tq٩qY{��7�vh�H?Յ�C���S�I��c���ϻ
[~U{�U!�#��;�L%���/�E��Ѣ������EC�I���w�����2�*�:��F(�*�]���M�S@m.�O��)̐�.xEC��5y�9h�t�&N{<_���V`�rw:{���Lp/u��47$"��.;� ���<�wў �4ċ�JǸ �ُ;�!�%�߯�[��v�&���� &a�p��^����'��|R�W�Y��\l:w�]�?O_c��m�=�~���[1�E����3�:��5��ʶ�l�:K°Ĕ��d�L&���W�͆U�vo���M�&b? �zzE=�v��**�"+��g�]T!<��n�Q��y����$��s�[�h�E��.F@5d��������0�f?�Ӳ?���e�0��K��0��B^�b+:��f��ejR�V�\�������j��ӸA`��D��L�|p	�^�g,�����/��[$�#�Cߔ��hj=>��K5C���H�
D~�-���-��9�E''���;8	F������o�E1 �"i)Nkp2��(2R1lA"��U���&���V��e����E���\�������H*��r�CY�?R���g@�����?^�,��΀�N�6�:�I���7����F�m����;&_~&����������b.����f�8y���ǈ9��
����S*DV��7����� ���8���|�M%J���6}�T`H����d��p����i~��߁9��)��g��	V0�Z=0V`Q���.6���� 3�>ը��,ƽ�����U�ػq��xe+�&����Ǧ=�R+��e`����*�z���~�*H�޹�I��0P�U�Eu�D`��tf�a��タ�kb�-����r�p��{�}�_=D��R@4��ƴ���	DD�9jҨVD�y�-4����9Q�11��P����Z���޻jSA-fbɬ�]"H���/���5���t���� $$�%��"�*v4Z����'ɹ�"��c� �8/�?)-��c�Y9-�����	N�i���ƽ���͔=|�u@w�b����i{�С�?] ����8�����[�i|M
�~	�CZ�*�x���k��3-�r��k�)=�#��p6W9;BdS
(*D���m�;���h�̔�YN����m�w�"S'���3��_`����cIdl�(nw��(z����0JW��}"
7?Jc��q�D��Ir�¯�a�m�e�n��ٓe4ն�C�����&ZG��}<P�εR�h�Y�<m
Z㻤"�Pֵ�ⱬ9Q�KGYDǰ��z郸�35n~Țzs��8|Ik��q�H�)�t�"�k�悤ꤩ0�ş�~���4ի�*�}��=ɉ��Q1������:4���JW�aj�s�J�\qրt9y�Y�M�6_�U5cK��=td@���px�X��F%~&�j�b�t -�썃���<����I�]twƂ�1���f�:�S�H"�! U_�������6�K�H���M#�~�6<yتq>G!FY��ؑ��Yr>�P�oҲoZ_n�5�ޠ�~��{%U����2ΐa�N����W+t3e_gxl�s���/Q�>���e����`�DtD��Q�LcIL=C} ���t �3��
�Q��
z'��۹g�w�=	c�������y0�t�J���O�5��B��~��lj�:��Tʝ�� ���G�Y��S�/�Dt�V�|��=}+���
����A���3vUՄ�O�G�|��x\��c:{^�Zf�F�4t�v�3r���W|��~<d�G�?r.���>�u�DMQfI�iVd{��qI�!0(�I���]�f���vX��p��]��9z�]�q2�K�ǹ܎)ˀ���	�1gEP�0��e�l�#.��5�|�@R��_o$F�!�������A��1�`�����<�sL�t�ǆ펭�.�_�����|X
%�o|�|Af�0�R�	~�™����}�]C��d9>Z��N��S�Ʉ�(,� ���q�q�&�,$�Ww�o���U��"�R����TZi^�lO���QZξ�%x�QR���܊���6�@wf2|�uI�h�OYu�dqn�Q��S��Q�6J��R�:��TR��E���*N�A��	�I�[������5~�%�#�#��Lm~�B�L�4w_/CD����Jo��3q�>	��}���ڟ�-��|��(N�kW�ZկeY�s2�8?xD�-i<���*�s:�IF� �I淅��H��h{K@s!�B���IT��T�M+�-��N�E����I�Һ�۠.b���l�<�� sP�eS���j{�?hH��=i&+�S5�
(����Ul�V<�Qn&̷m�ˀXw�ϵ)��~Kocť�ǐ=i4�̈́�E���v�ɔ���䫝����J��h��x������ﲀ�����]
D��wP5���LO�%Z�e��T��Zg��d��k��ʄ*0K�s�!Š$�΢$��)�3�G�K�V��*e7��A�t�P�G�}$�!��eU�rUfZ�Zz\�� �/����L��Ij=#U,B�ςScY3$����a��4�@(�y0sg�b�}�G�����:�w�q8x�/�沓���hT�C��6����w�#j�� pC�?�Q�Wacx*���J����Hgn1D�!�Ĺ�N(�y,�+y�x�"Lܿt���
��3�Kbqik%�`Kh�f�~Bb*��f��\�_Tw�d�lQ�hk4F{$��]. p}�Xٟ�{8�����#)�1�<�Ub M��r	u4���Zs��M9�;>���ܑ������[I�ⓥ�Y�q%�����ku����c&�+l#���������p¶��
]�l��}��Ģ��j��[�0������q����g�>�����K��g�f��M"!���ϥ�s����^}��/O�o��}��v��'��7�U�T��	�}��;^-�I�����F�gMvgĪ5� �<B9\C�~r��2�*��\1�����ߥ�do]fei�Y*�(������d��F�X�*A��������#��mu��ؑA
T�F6�gY�������~�	9!�L�������/���E.~W�l�
�.7�ѩ��L�X�����T}N���.��O�Ab�����#�lԀ