��/  �^���H��r��l&��O��,w���iE�d���S�d����ˆ9�{��$������5En8�k���
��1qG1��#�:?r���^��Є8+Js{2]���
a����}X~�s�n��ab�"%zT\���_�\ �D/x'�䈹�Y�W��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n�W��ߌN��5=�8�:N|���gp�P�ظ��U��)�& g�J����[��kxO{F� �N�2���~��y��Fe�R���n�F���4���P�P:�ܩ!�{�ud;�魖�c��B
dM���u;�w�C�$�-�����Z5�9���HR�t��S<ʐ�t��<>.��F#
�S�N�|Q��v����P��F�[n�jnva�P@�&�߾�t�����gË�3��jr�A���B@���.�I��~asDs\|+N�_��B?������>~>&h`��+v�Si��HNN!�j��p̒�y'�ľ)S�IL����+�� ��U�[#-��b��J� �e]�o��8���:�Ǡ���'���{�.i�0Z4�-Y��T� ��ƻ�����{�sd������x,-�r#�.����	�S��a��#�D��1	>����tvm)a7*�?�:d��d��8s���c0ZQ��!�$~,�������Ǜ=Z�F�>��3�YHt&��4Al�����cYH��hMs�m��	M�hC ���+�V�� �~��6��0�E
9o���!�
_ί���7+Ō�J�+v~ �����tmg��&rCI�n钌�ʶt!�G]D���1E�Z�u��BAOw��[t��!���mK�����"��{ �nJ8;���A�J���^t5���Y�)"��V��r�49v�I�uT��Pr����X��	b��y����������D''p1Ow��Y�{��t�hY�H�8���gwK|�s��tT�f��}��5Lw�d�Q�␯�.�H���p\w.I����mnp���S��}�cռE��EU%֚�qZCn��A	����t��}���/r:),L�T1y�	�2@(Oz�ёl�a���S���"q��l��y��S1`d��j%�M-�����'��F����Ɓ����v�^�G�[�0�y��y*J���T�ң\������k��|E�M���Oyk�hQW�14˜��3�����K�㠧���Қͦ"I*[�9ʊv򑆩�U��^0Xzi�nd�������b��j�A�5��p�VNJA��"���C��=ty3�-q����b���o�[��l�b��[����Lo	��wg�XD��@�$�+dYl�_�pP�y��2�`�}��\�C��
sk*�-W]/��U��u.?a���T��S	��ֲ�8(�A�=v��·�fe���oQ�ev� K����� Y'i�l~���2+䬼9t1�e���\+-v &}f�u�� �z�Џл�/?�F,�;H�y���X͒v?׀�QpuP�,X0j�y�g]�L�E/$d�f�F����DШEm*?�I"��o�ƙ��4$?N��m�E����4dif�> e͇�����%pOlY̅��_O-����8�vb��n���3s�e�4�ƲӶ�'\j��J<�R�K�47�j��(��������3���K�IX�@徊Pw��w�>���}Gϴ=��\Q�c�^�L�$�Dp"w=��5�M�������d�}���hK��'����<"Y�Jw����!H�E�?TX�9x��i�W��0��"�F��;���R�s��Y�9D�S�&Y��S���jS�bSʏ��sW�ؒ�f���k���1��-���J-wJiWsm !��4ꫠ?��q�7p��!�����⡗:ɜ��+���9I�%�8>V��K&�{���-�Xwu�c&����qWx�iL"`\2�Ŭme��>��HP�W���`>٥�R�<�n�oC�+�-�� rYfzm5sx�����Q�=��f_x{�^ph��mA!4Z�j�x!���MSgc�St+a:���z��J�ѫ�r���i�bL�\��x\.	���|�bKp��P5��B�R�
���]�4?��W�ר)���"�+� �an��8[C�RG�|GeĴ�(M�&6�_T T��1�]�dF���-q5 y�nv�
�-<R8�~�@�ooOF��Ş���H0���q�O~��N(�K:㬨K� Y�e@�:I�!�����#����%m<����'/4C�H�o,-7$�s49 f����X���='��Sݽ3��c��V��%"*�\�\���"Un0�þ�@^��ǲ��|�K�hxEl���7�ꃴ$f�@�y�4�'�UJ��{2{%@z0��gvW.�t�����@���tQ�Ĩ�x��QT�V̏z���S����Ō"6a=�S�[?���3����G�+x�k8i:�`q1(L 3��a����Yعik���ڟ��>!V�M�f�b#ʐ{č�|�9N/&dp�.j����bЦ�]�0����_��=WR1h����[E�EW~�Ypy#��j�Iit�YL,�>�ޚ�u4�ɍ>�_�}[����<���M#r�^޲���m!��pGe,V��D�a!��n�!e2�]�7�I���9�M瑽����U�˷�ǒj�<�b�z�vb�d��h� ����ҟ�#·��'�4	�K�jVF�߃a�D��'b7����9J���]���G.ևZB�g��M1�0�;�'�x&�hs�4.��J�H6R��`Џ���QO�[���&g�"��{���=	�:�$��2�'�6��(�PH�ڽ�A�L�[͓k�̺(���Ȕ@��լ�Ч߫�𧣫��q�c*��Pw��J�JM%g �=T�n�Sqa����J����^ �4�E�` �1��/`"���:a��w/���0�H��%�w��xC�������pĚ���F�<������f`f��6K��T�����j�R�MG���W��3�v}_�*�:|O����a�)]�Αݽە��庁֬/�β���"9B�B�,~��R<���V��F�cS�k?�uT-dQ�J��f�3!m�[�FJ�]��ߟ?�hj���I���<�`�h�d�&<� D�!4��c�+)���q�{��	hs���+神"c&����7�
�X3�h�gNz.+;!,b� %
�s��%n���sDFf���}�=�[��OƖ�3�T��~�v<C��Y<�GN��.R��8|�L+�.K��J����U3�V�4��k!���@�98�R[��߸��x�,�x�G�G��Bfn�S��9<$=?ʁ�
�_���\��o��]D~��ZJ��W�z :�^��9�s>�3��-���đo���:�0$YPґ�=V�C��\ݠ��OA?2�����.9�L܊f�tWpri8� PB.�Mq�E��s}k���������F!�??� ���{
F `͔��Z0� <4z��0�?ח��#�7N�gNwCxÈ���7
0`�����0W�N�l�3f�ofù�Q�l�f��=Z���Ǐ�jkb�')�';�8~Kw&;]��)�f�-���.m��3K��_��U�t"�N���vCb�
W��{&�oi�_��V�X�(H�-Ŵ��p���m��9,��ڦ>��Y����,'�Y��[�i��;��)G�+r`/�*�8P�/�v��1@O��#n0�r�G��=��j�B��B�"A��>�NM��]840zy쌓m���Tk�V�KŎQG��]����,ì,_��䶉�6�l���0�b�>���S����O̡{����� ���Q���t֕�}��8)�:�	�P�p|$ׇF[>^Wޫ�����P��?���qZ	�cR,k]d*��@e�gGE�טw��\u+�O��g|�SFhԽ+>�`�Ǫ`_���($��߇b�%�9�F�/f�P/{�g� �bB�8x���qI~��?�[��B�B�0�n?����%Ӎs��