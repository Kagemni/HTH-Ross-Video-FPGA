��/  �}�Gl�cV���â<��������qx��Κ	˅���gD��0��7�*پ,��)���R>탳.�Y3�_5�6�t��`V�e˔��0�̛����h0)L��	�W��؈/DP+Ak6yfd�%E����u9�摚��8g��,�ޟ�p�Q��eгC�Vq�|����D�LDz� _�K2��({�ya�Ko��5�-`FQ��r9������
�r�Ȧa�z�W��T� %��֦�8��G�BsqAױ����[CR�ʜ�K�|m��#R#9��G�Zx�g���g,;���D�;I�M��no��h�w "㧇d���?��1�����)�I��Sc=Za7`C���ړ�(�9Aa�ghB�E�bYQz��
:s�'Ұ_�3�튽��(q�)�t�^���Z����*Ƃ�~�D�y����Z#%`#�r�V8�$�Bh7�n�r�}�#��e�D��ob�|�����E�\i����M��/����Ǝ�G���s��x�kB�,�?��������~�VSn�9��no��h� �7T�AE�l�����~��jV������J����f:{���pnD�l�7y{��:p�U�#��u�W����ПC���ҭ��c�����'����\L�"�M8�9m���"�N�;��*[�L#����qj'�fʲ��̼������_ddE"�kR�b>t�v(~�$8H;
�����f���l�a�|	3���{�+�?U��w��xS�U����r���T���7��#�s����峝!�R���4p�$�зi�;���d=��F;���%�y��iB��Y�܋EI��p�����FQB�X��)�r��!��V���z9���չ���Jf�+4����AR�方D�	3._�zww�G����1W�2>�ai_wN�?�PE<CܯZ�t՗+O'锦����Է�f��k!ϫ \���;
���1��gfBNo6B,o����uʌV6���Y^����l�`�J����f��K#��Fo��'�N�z�G�3��GC�8Js�`z}�n��/�9Oi�5ϋ�T�cP�"I�m�pC����ekm��hE
��tk���(�&�� ~���k!S%.�Co��&j� ���J���Ԯ�%�db��4$Rk`YGJ*�pgClQ/.X�����R�����mQ\�b� U�T����[{��U!G�d�T�@ ��+iȿ�������jh���ip	��+������T%M�B\#>��}�GC��%yH4��!����"Ui�֯���+�Y�D!c��v)s�@ ���i��%|�F������E��8r�$�����·A7ܖ��]�o�!�G��W�RF�}EF_� 5��Gӱ�����0��%��{r���7ՠ�
l9*9�iX���=�J��I�r��]��9�G��
������^�?�E������Z�с�K%�\���QpK4"*ڢ^�6�c�	�)����U�w���
L��w�����E<��?/�nmHZT�g���dU����e[v2.�z�x�e=�t
EP���B���$��Õ��=������E3��NX�_�*��g�a;0��<� �G�ۛ3k8b'f��de��A�����o4���+�Ĥ1w0�ɔ����C,�Ӫ�<S�s�j֠u(?te�Zu;���9Ҵ���C%��6/��~�Vs�"�)0R�:��2􃌏��?��E�zT|�� Z�2��G�Y�p�^�:�}P `�����$�OO��K&��L��/��?C�}!{R�4v�3K� ���]f`� � �TyR�Uq�z����	&��7 z�b�f/�r7X�fXt��/GIֺ���;(	���J#�;��%���2��[�d�OR�ʖ�¬��(�pN}�m��P��G�3l�8�N�?\y�D���%�'��qԴ��#�\I�a<�xbN�� ��s�Cm�D�->�Fzڡ�%���� +i���+�{NΘ����rLb���iqt�����q�Gj{ϻ�+0�1��l�Ԃ�0���Y�X�l_�v*�ϳ�t ]��9{?�B]3Z���Hw��?#S)yD�������6��<2|�
��Β�.L�r�f8 �q��	E�N�~�}��P�3�C�%��]�8Tj@��
�A[]�H�cB��ˇ�!�zI�炁����"�<ьUR�Lv����ʏ�6IJ>�| ���A������ڃr6�?a3Q�"�@��K!<�.0�}1���U>�׎Vi�?V�F nU
�QB���\4�U!��j����8ShЅ;r�؊s0ǈ;	�@�F?�| �Lg���,��=��ƒU�h�W�H`��.71lD_;�͘��,�7�+J���ds�Wu���i ���kة��g �**�m5+E@��<<�0f�o
n����:��*Ǽ���0h.�~�.Z��h�Wɲ��Vz*��������/���l��J��+P��*��o2_�י2,P��1�T�U�ܨK1]��
P��@��'#������n��"QKPQ�m�� �b�F��ߊ�� �rCD�Z������	��4h���?B/r��i���ܦ�|��s޲��\���Z���2vL#��;?:+8%����{�$X���S;O}]�@м!����6�`�ɸ�(�֤CZ��_�V�:I�g����Q�<=��g1���#�Ǵq��] ��WY��r��ȇ���8LIb�H�
`oƻW���n�W�l?�q�[����ݽ��φ;�����ұ͂/@����*�����A ���| �5�	�d�$ �9,��ލ.�'�솜�%�D��t�ɻ�_��R�<h��#�h�;`�D���$��~#�HAqbf��;ч��j���.NgK�`�I�ʞKa��¡e~�9?В�;�&�j�u��_��t���ǡ����<	��Y"r�(TO��28=���<8+�(;�������2��{�_
Sk޺)���a�ʞ�ɶ���3 ��>�(�=�:�ē��l����W���˿n�2�v
���QK.�s��sh��1�E]�UCV�`��������@��_��挤iR`�$�њK�Ģ�7���z��r��ъ���2��>�n���jkNԌ �
'���6tG�[�����S-7g��J,�3���v&[����G�e$OOP�Ց��)�ŜZ���p������*�l�|�d�a�6v�a��3������zcq����G?�*,pL��DԎ@٧���� �-�{I�v�^#���P�TdI��}�HM�|����� �F��V@�MDnT8���;��ҸE�>�|�t�D�B���V�$������XWUϚ�W�i{1��%�Q����d9\]h�h���)���q�]ρ�K�Pn��ۮ�G��aR�mo��[ ׻�i�So�:��E䀤��<6��کm�96H���m1+�~`��HrvŞ^�a��e����I}���rQ�1��B���1�[���[�{��&u����ԘUX�2��d̃�ǄO��6�P{���S���[IF(t���}I��6��]t�÷�ƪa������q� (��Z��o��\�F��e�a�F�ޢ^ܨG��y)�� �Bm�a���Y4!}c���4//Ȼ�{��xk)��'oǁ��.{�H\��b����d������2V��B�;� w��gZs)��暢�TAi�-?׺������a�R�L=Q�ՍL3�_��?�^�x�5eYtα��F�]��:���y��K `P��!T!q�����K�� �q]1YGFxl�}-��=#c��fg�s.`�/
����W��<�i� � ���17��#E%��Y��P��+s��p!Z�JE9}�N#���\��8:|�T��vA�*p~�c�A,�e�y�dPe��Ct(�=I����J��lƮ���Z��z��k
��E)F�N�e�θ���K�d6�Fδ�?o�&g�fc�5���V$ƫ�N�
#�&�����%G�T���/B^�z��̂*?ݝ�q�g�ӝ��^ȣbLI�*������