��/  ��)�����p.o��;5��}UIO�1j�āw�xN$��4���8��S��F�7�];Dn%޻�s�A'��@�����j��$���ƶ�E&@iG�����:��`�h?�����k�Kxy5m�-m��W�zyyrڜ�-/;��޼ݕ8�9s[���kWI��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n��=��W����9�NCvZ�gN�%#jg�5����u874-6��*5.-PT�^"�R�N�/�n�|e�ßs���=� ��Ӫ���b�_[���97�g\u���6�ȭ��e+��ȩN�\tw�T����n���X���:�f���;�^v>�
��#9��歨9�<�Z�;b�%g�=jC�͢*˼hb�|c��ƒ
G�ߚ)���,8bt�ަRP�}��C�]�_�㫛�'��"S#�e|
��*$!�����5�|�kYJ���j(���I,7X�ʁp<5w��e���k��HK���#k+��a�5�a����f�Q/�N�T���D5�Q9�Ka�^���-&<8 ��BS�	Ӟ+7cދP,&��I�E>�]v{v���}�rO� o^M��t�7T
)[��~�H�Y-|{�tBA x�� �R�.�5y�a�@���mi�=�aP�+�""Uf%û��oj��e�2?f�a�;�T���X����.��7�K���-E��u$Ϫ��B��3�B�,RrKv�[	ק�wh�����&��*hZ�]��t�����^L�^o��S:���_?�f*���5��$sg�ƚUs+��0u���)ΐ�^��v
����>Z(���99��X	C)�i�8ߢ�ثfd��2�L�F�^~I�e��'���=����������te�.�\�hO��㋌�n�vh��b%�p��r�����T�2�3��r'�Q��u���_��*�~�������QrB7MD�(t�� ����+{���;�0�������Jx�2-��L�NyDTs��
y0��l���t\�h� Ӡ򏩳G�+	��sD����w�p@�&Z<0���1�D}c���?���/�GPH� #���}  ���y4Rγf�#�r)zt�m���\7�&ųy�o޻�q�t�sb��ڄsm1T E1�:K��~���S���U���Q<	�v=6��;p�+��[����f��Tƶ �iG�e�DM��c� ���v�{��&������ဘ�*�9�RW�$�`�1�h)^1o')���u�7z.�+/N*u{Ŋ�������هş5L��ic��]�7����*+�[�Ze7ߝ�P�Q=^x��=g�7��a%�~�iG��+�Y/���t"�Dʍ���Q��ϋ�����} �f�3��|߃G-�VD���^��{��t˿�P��\�T��(��#v@{n3p��!_$-����1�IT���6�
)'� 	��~*�8B�H��i�]���z��">�C�����ߞ��h�I{m�~�tx3�N��kSJ/m��ɉ����%�D82���۝J��JOS>�)������e��&�گcV�$��%8JE�?�ch=$}�}��+�VH��Q�F�zJz����814� P/9���}���R�42��FUq�HYp���⣘��Hf��� B��?�_%Px?�Ԃ��4�^p��ߜ�>kŕ*�<Mo~g��mᮤ����&��/�XU,�%ޯ��5qV+��D]�з�/�KaN�o�r�f(t� ���ǭ �~�Fi/�V6>���WE�ݙ��6K��6���%��Ԫ�S2��K�?�9��_�����ա'~F�k#���i:��j����W�a�)����s�H�/�ڒ�9�m�oG;*1)�<���=�0��P4��{��@��Ʃ�F����X��a\䔰\-6��R���,e��,���z|�<EeH��i��6����[��6���8JÇEl���� A/y{?U�V�F��������g��S��y�����Y�)g�dmo�)�3ۼ��b�S��f�פ�G:E�8�%�E���Ѕ|����ߊ�u�,�/��iĂ�6E�}���?I�l��h���B�bl��{�7���ag��@$�-�,�ߍ���R Ï S��Dʜ�䱊�N�:Dn���h��CN�Ur�F������k���]�'1�n�6��/���|C�s)��yѤ���0䘢.�&��zSE�_n�����2����j���-Yۦ��	ML��g�!h��t:����
��:�����x�~� E!��*�
�*�؄X���Fc4�O�kRV�������!��윿"\m��Yp��wi1DH�����)Gʲ���k�n/K������RvT8a3�c�������>�IT.������k�X#���L��֏S=�<qay���@��j�]�j��
�#�)R�q�)����-��!=�'f������s�cǸ_����2W��"��quJ�.�wД=����r�n��4����vr����@	��Go�8Y����h[�!�ci�ġG����꧖�t#�_�<���K\��+�>��@.�Yp����
�t���b~Ϝk�`7�+�q�"��h�u<�:䖬h�Bm-}N)H[����5L'R��G�����rS�w�I���;*r&��` t���J��{��v��L�.�;��b^K�^��M����������2�X�+�,�����U0��$O�7h�����"a.�z>%Gב	-})�mzN�%�'�I�����낈&܏շMk��U�K�������� �B��O�]P�i蚧�%��s����ܴ1����
�(	V�b.N�'`�����Ù��� Us�E1G���N��e�e9��pv��i�ȞQ���{�j�����3f�A�ӣ��K��fQ��G[gW�o[��Ag*w.X�����z�|I.�Q&�#W0}�m�5(� �y1��q�C%�/�A��jnTBL��d�q{nǘ$5���b�G\Ms(y��{�LIjI=K�.�h���8���p_=Cuڔ���bPI
���n�/�7j���Dc�Ysq-�Y��7������q��V�w��&��������~��x��y��Ĳ�l@����Z���f�U��8��?3&�Q?
ݝ�P���>17��y��I�}S���Q�c{�+`��BD���;�Dʪ�K����� ����fYv������E6%�@��⸳K-���Ջ���c���	�wjj`%Tƻ��ť��4[Ym>�lx�Ǖ���p:f�������d��=�����3~EK���Pzw��f�m.���[��mn9��@�f�XLZ4{J�oц�e@��A#�H���Ƈ!$�H�����	g�;@�x���Xk���}s/g�\u��6G{v|���Kd@��3�
l��a0�9�b�Zh8���ޛ>�7-��r��T�\Ѝ3s������0: .�g�u	������O8���L�3�PՒ������@�����p�P�a�������E�yU�!@�?�d�u�W;����q��#������؉{������vO��3��:�i���&fԠ������9�N�N.��$�p�/Hna˭�;���=�>�P<Ι������~z�\;?cwN�ub�����0����l��M�~�?����>�~��f��]a+(��'���O�>^u������I��k�������[�/i���4�����p8�2P���^5ς��[�%#�v�N��Q^��{a�9D�4�d�	8���V�W aM�Q�o���dذ66Mj&��
��%�1�ݲ%�@���J+������
�UYaC�#\ �$� ��? ���s.�aѾ���]���a�:�9�y�N�s�S��׷�l�X~d@��q�C9 ^�N�U��=�l���J�7��-�8����r�fhc��{�<3M�Yů�O�'�6"�2ɵ�HFa3����z��:%�=�'ݶ�%P=�IT;3��Uz ��5zPd���Բ�y��+����|��T�w�N���k�@��=?��@~J�ͩPW��l;��!�l7��[�����=
e���odx���1���� aQ&�?�W��CD^zbǒb�[�i
��$�frT�a�`�0�|M��<�����*�����k�g��XH�q�$�4z����Ћ����PX�d?nU"��hP������}�}uL�<T�FU