��/  �I1�J���%.���z�m�l�����w	jݺڪ�Zp�n/3�&��)&����2M�1h;1��xz��~(��qH�ZÓ�N��� L��?td���UC�G3�������Z�+Sr�)��@�X�$Ͳ\�����M��>�Z��ۋ��y<����4^��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n��:>7ߎ��Ғa��H�Ɯyї^sXz�1>l��^OɧF�e\p��.�Բ�O�mVZY�5F� �~#�:�Mܸ���k��6i��������u�vpZM�r��|�D�!����<�&Dn��lT���$�E^
��֥mRR��G�ѿ��D�VI��5#:"�*( Td�Oy_�N҃�&��B>L�~�e%bR�-[�܆�o�)���l/��7	������w�9�gA�p���ԙs������N���Y�x�H_�4�T��ה�#{v�������Sh��/%-�|~�]wz��Ux�_Z��;��gM�E���j��\h|U8�������\Hu�CP��ʦ��7=y#�Z��Ϙ!<����Fg�4LQOm��R����%�R�����t��?�7T��=yk�oj����?m%����q(=�xo4f�K�Ǩ��Ch���<8����{����K���ހ�WW��t#��}o6�	d�]�{�%݌:�s5?�K/��\�x� ,p�3j+{p�P�w�<Z�u�쌐3��gzӝ�nt�8�-�ޔ�W�������T\��,N�v���Bͮ=�����+W6��$߳1�P�}(ѼL�Xi�q����Y��[Ӏ�ML!��G�ct�J^R6!��S��"x�4���q5� �M޹U���Q>��>��ǍU?�L4f�J��^�{z�$Ĥ�nPN|�jVM���gc�wV!N+����(��]�Q�tj�1^��Z��_��1JOx�rJ��*T�~�f���,�zCܵ�=�Ir�^�$�(��;~4�z,��o�
�ËM�n�C�|��O㤌�e��R�1�u�Eˤ��tL?>B|(��a'ƨt�1�����|��҈�66��zfc���=K9�~�-��ƒ9Ż�)�;��s]���iN���9�V r/t����5ح�H.�2:D�Ec�y wD�uG���sߊ=����Q_�Εu�L=����I�kR�<�L��A	Q�U?BD���3x$�~���SU�f��|���=V#c��%B�I�����b_&t���g���ij������%?�1eX�\;3�Y����[պX�P�=n��K|�5[qɇ���(]�k���g�������T��B,{	��8�"nT�"���5ߐ�O_��y�z���թ�.�Y˚�<����n�:�3��}�,����ts��O8``�*^���i�̭�b��7��;�C���9�i��hJ�C�$jܕP����n�*-�8Čm�4'�]kq5D�$��>�s�8����?E�����o��Cd�yg7�qaN�hӡ����{CDu)��-@�������ۿ��۩�C�˜�����"ِK��"D��"��m��{�͎�;�d�a�M/ʷ��k����)�Agq����K�$��lk�J�����B\[EQN�sC��E��zz�瘪-M�W��dK��9�,�].�J�e��j`$W�[����[ƭ���o�/p/t���-u���3�;�Y�&�1.�C���k���Jv��+re��6�:����!e��xq�c�/�[nCުP��G/ŠX)~�~,�|+��j���L�{�:��>=Oa�Ev��᳐�[c.rT��[��6�l(�=�{p���Ei}���?������K�R������(�h�5���<ר��wQ���_\�B(�*�jҜ�xL��XX\�X�F��F���%L_B�"Q����ѝ��GP��2 �Y��q�[l����/$�������KY�ǋ���k`����Y���g:�a�/�O[�Epj /����X*���I��㟣S{yzo���N�k�J��m	ŌF� �L|��$���⮒Pd����r���oI���*h���"�񍭉Z�L��g]ha���i�fI�ڶ�c��7	�T/9n|2���J��W/��|�Y�BnN�8�d��I��w�h�0x7���Y�/.Sã!op&�1M���ɂzۍ��m�
��$�I�kG]u�/��*v*��-��/�B
Y@'��h��y&���#W��s��󏕁с�Zi�|���W�J�=��Z5��K���t/��j$���z0��w�	����U��maF�=�1�t����A����#��&�K��!�,�(�;%W���?@4���-�Se��̻�#y8ȕ~Z���!P���&�:�U�UP�l� ����8X�]��Kz������r�h�1Fq�{,���:�XAsMo�y���S��m��5�y^g1�0Z=Z���@�R�д�g�B���<�GO�����|:jp�@9��>%߂�S2d�$��0�92�
-�5�<"H#ń���|�s���v�^<zGI��*O�D��u��an����f�m*�#�����p�ji�Ta�����Ze�f����G�m���m�̞.���>�$k�༬-�h�~��a99��_��{�e�욮mn���Q���,!1)
� �
 �-�6B���0RL�����x��d��VO��\���\���Ȼ�k���ro׾M%b~s��{x"a���t_vXw|�A�|I�`p������{wUV���(�f�5���N���?G�[�n� l9�)��5�v�=A��Ac��#�bĎ27>Cs)�Bb�
���a��n��|��uY��!�-���I�`�P`p^jJ�(�3��<��_�ߎ��"�9���ƿ!�ͩ2��ʾi�+LHy���Ĥ ����N��ʹ�!)�
�����U�ޙ\�p͗(��Z���R�!bW�>b%Cl�';�@�j�����5�ߔ;�2l�n띢��p&��zLe~�]8�m^� .6���W�8�j}������[��L�v�#aPD��"3b�.��R���� C��J�p�˜),T*���!�o��,�c��	��xN;f����T�Y��
��bAPX^A�����.���_����#3a�S(?�^�=��݁��u�W�Lw���`fPG+�����ݡS�)�Z�JrSmJ��R�qp��q�	��?E��Yv�A�~eH-5G��Ap�/ �f޻Z���$�ThK�#���U�u$�K��ӓ�x��f