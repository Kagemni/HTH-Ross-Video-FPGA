��/  i�`��,��j#o��:<}]j�9j�T��lo[���R��	�8S(/V�:����/RMym�E��ǀC�2����!�"
���Y�7Ad�h����7� �5J��U$'I�	/��)Vf�`��ڣ���攑Ł��(���9*	��<��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n����D3ӡ���p"�pM�x �GIc�W�	� ��S�w��Jƙ���� 	+<1Y��O��1�bh����Q��"��dy԰�|j-���F}+g�`|��Ѱ�}�؀L6!鳚�}�؋���,��>���G��kw��Ζ^�W&��Y�3��T�)*���\��@6N�r��D��L1�,׏E_�hk��l��5�G����ݖ���ݘ�>�F��;��*;��Rs��;#�6KlLŉ����C�^�0V^�錳Ӭ���b�\~&ZU��2�tz-��^�k)0׉& 9���P&4����.�8��)]����Xl��,˚��)H��|�B���)����f.+�������9���a���e�x����Rlځ�u�[2��a��8j�tV��m5��p���]��|z�,+�N����l423�t��-Qf2bB�O|�/!s�´�E�0%������<1�U7`).�����|��|��v�H`g+��WN�b��o���mI2��^�	�V��!zc$�����%5�WKҗ�i�E�ٞ���}SR���YҠ���)t��&����t|4B�zAQS�)��3����1p��P�&*u1.V~���{�՝g0?����ݗ�0��eHMޤ�K�����#�	�Kl	#5O>�"c`��`�6d���2wj�W�A���F�xʭ��Dʉ5
�hy�e7��~����a'�9�zx%���Eo���z�u�5�?��JHT�y�04��<:��E.� }��QG*&��? v*')NI�=����#�^aFF�\�Ư'_0aF/�R�-z��[�r���P_//����re8S]���?�GA6�{���cV����]U�T�S��@�(V��8[y�䱪*�|G�ƭJXm�"�	�g���>���}��M
�	F�[_�U��0���l��
���JM�ٜHp��g�	��ué�>˦�ƽ��3갶ۋ[ F��eR[*���w?��b��e$��U�6=�~�Ee�Gg���V�*!�wN5d�؈�-��+ql`Ps���_U���Q�wP(f�x��WӲƁ�Ý�lv2#��F�I��W���W�����>�L����T�oE�,���q�Q�|����n������j�ވDҁb���Y����O������P� ݉��&��A�]��^�Cv�l|����CqѮ����1����ۃ�N���I.��A��; ���
A�̜h�s���sP2|���6�VR ��NdǇ�d��&��"+BUI���{=�d&��0{����!�Vϛ|H���Kcx��:�#g>���2<�6�u�H�ND���]��i!�zhD�����M�z׿�]!�X}6�v���s�~Ē�M�w�|�[.yq���?p��_v�W�à�C�s ��Ձ���H����
�Zc5|��Q�mu�RAfĜ`�XcW`��v9`?����,UiD��ua�ܟ !Z����?t2��r����Ȣ������iE��<�����Gv�e�Pq����i�>���:	�5�P�<�q�I���1���"?�6�����#��I�&⤁����2P�Ǟ�t�zE�J��q���&	�0��En.e���o��I�j�+e�SӾfB�m��gN�]���QC��/4��ܲ/L��_�[K��}�X�)ఠC�ۊ�kE� ]�!�լ�c
����b�i�b�F�&��>�݉Z�/�j���~�(%��z�3�Xƅ'k�޶���7�����Q}�9Ep�l��[�_d�S�/��a&��Ŋ�bz}����
N��A}	ր�А���c%Ll+3A(���}�#J��C%�g�zסv=��Q���[�Iy�nʶ�@�a���ļX�ͫ͢���B��u[k��#��jb����k�
x�{u�;��RYaP7Y�|h��ea��\��n�i�<ڛ�[�"o����R{��\�R�,�f]]�؟�(��]�L@����I扈YN�N�G�*<g�_-e�K�KH�ʏ8vZe��=3��Q���vG�ͳ������A��D�O�P �q"M�QD*�(p>�
�DQ��G�4��k�Y�pt#�I@k�=��r0ŵ�Ǥ��"��m4|��sHf�]˙f�d:��̠o:�X��o18�2�;�Wi��(�%	Tm��D[��P4���<C����Zn3��Dd���%��@Lh�1���%�%{�٨Ò|���P$4Um�G���7L$&U�by}��9�A��+�v�%|UYȾ�o&K/��5��%�T��0���Ł�K\BS��l�'</��N�4��X� |��'�X�8
o�gD�
��%�����Y2���
�-:2�,��CVc��¸X��fWye�u2���k�mRXX�ß嫝��@_�x2��W%��/�M�v�CD������Ub��^��}BAQ��5N(1ޝ���a'�S��`������JLH���8�J�"�1k-D�E;ۀ�ؐr��#:�q����v �����*]��1v�W���n� 8sS�d�"΍s��U��g���� �0�|ؾcjze�>���B�;>m!���B���-?������ƢW�׾��~w[P	��CWհ*�h(+O���
N�w켰���1��Q�Җ���+�)}�\�Yb�A�fՃ��)���Ҷ�P~��Y˓ڋNU�j-��H�<x"�0����0�D�s�����)��rS�9��Ȓ��׀�
�Q��6ʜ�jױF/#E60��e/���b�n�fbqע�,bCt��l�)��"չ�Ɲ5�=�df_���آ�X��\���bUt���}�����5��"�����[�-���bfZ�qݥ{�^}�3v��4��q�ζय़�8�XXki��4xn"����S�
Dc��{r�V=%�s���ȗKMZM~��E� �*U6(q�>�S���T�ь��]'�7�I3�`o�Ӭ'B�gn��/(u�ڍ��7�Mф�I��j��,>ryI��0C�]����;������]���3б��;8B�tu�5Y�	�Vs�G[^�L^�cv*� ;FpN<���m�rڏ��{%?r���Y1F��0�0̩���7q3��O5/��%r��m�^.�	|�M�������)�t�Sf���S��xvd�4#�U�kH�k��p�V�(�&~o%_�5.q�\~?���חr�59������su��@+E2����a�����}08���RB�f�b���0t<�#Y�q[1Q�JLV�B
I����H���"��/i�bӐ�¢�Ȩ�P��p��A��q���᷎=���G��p�����S�ƞ�4��$"	S� i�ڢ����z�ގ�9��)5��ŪeR�@��ͭ�q:�=��4D�!J>ϷS|��W�V��:0��Ŵ�2�*O�W�`|v�m��17-t3~��U̵��O�J����Od�D�{� �Xo� 8��k�>��qU��2���`7�˨�Ͳ{*S��W�u�P^��n#Z?Uobg�1�@�%|f��K������F�|��%�o�)�d:iN�`���A�����(S�M[��KUu����th����m(FD_]o�tYj�h'��yJ;3��;uF�/�P�?�R��:U�K���������3�w�4 Ȫ����-��5P���(��՗RZ����;�,d���;}��>���O�~��JI+"i*�1�������N}GKo���3Su4Q�U�3�%�z�H���J�Ɖ�xw����4��J�o|[h�~�Nbe���[,�D,qm����p"��YgB�]���-J��u:􌤱rW �s��&A�&$ �̤��0x�W5��5)T��鞭,D�T!���z�+�p�b��
Ί%�J�[<���N��){�����)��ig)g��e�ǚAUR(����'y�߇���8z��h�=2|ǥ\���ߺ��o�I�O�|I��`s�su�/�H1ߪ��ey���H�wp��Q�O��hC����Z޶�L� �!vK���Zҷ�c�UUޭ_����I��F1=��K�8I�75���5�f�D$n���16{��+�?<�(9{����2 '��%�c0��#˖}�WMjE�Üc�!푪�y>��0���d��:@�͂�A'�Gpjɜ��чKj#�f(4+��*Ԗ��QԂL]�}�|���?8[D?$w��G[����Z�6Y֔`�`J԰܉���d����BrRGdǗ�!��͌)�n��a�$h_�����ń��A�`}�(:�GZ����<�6 c�1�cQ�Y�)���̕;ā%�qJ<��O��$�]}�lxQq�,d��N繇��Ŏ���Q�t�Ln���p�9������+4�Y~�bL�L2���^��B�����s���3�������ȪPz9��,�H��^Pd�Wߒ��<��JH���K8�4p�*�`�3���]��׫�'���e��>���߬c�̝0gV[7�6li���l�}�tH���r����́�VڛVE")�[W�'�ݖJ�I�ޗ�Y���}��Xb""�0@Ԓ*�<��a�ݨ�_їOZ?��Z8����Pc��8mɏ�
�z��4�vAY��n�$�0f�_o^GZ��R�<%�H�4Be	�f9����4q4��������/x��lvHܚu�?}P�f��P���?�zl�����2@&��#
�G�b8,ž��7��of��r>�T����A�c$Sei���	]hqub�-�_��o{z�~�#M,�M�r�ϗ	��ë���u���C��'Ǆ0j��K߆of�b�~P�����Lq�&îa"���'"uD��cG����դ�cm>��I�L��T�#��Mv��+���*���U�Ӣy҅�O�
hr��+.��1lU#������n9�"��#k��ߚ=7R�u�[�"w�!�T��66�zLl0�