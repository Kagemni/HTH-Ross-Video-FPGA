��/  �����d[�P�-�
d�*Zc��ۛ����X�\+�M�D,��6,Lsڥ6��c����L�N��7��4nX,-��v��C�����;����#l[~��0�� ǖe_�@z�8^�(��l��I R�j��|k���Z^V}=&Vl	�D�I5OIH�㠏��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n�||�p1��b<o0]�z��L�^6'
I�B��������"z�S���')y��oK�W�xZj� ����s[xl�a]e6A�΂�o%5���+w�7���s�G��( X32=��4h���3��k���$�ُf��V�(붲�� ��?��VJc`��Æ�tU�I�Q�+-y��H v@M���J�6�v���N7Ed����wT��������w|�u�%�q]��Eznf��sc�s�h<�E�@v��o��"R�U�z��Wu���3	���r'���k_�`d����}���
:/ؖG�'Ƙ����{�fl���W	F�M��=;�^���B�$���=���bj[%�����r�H�-ڇi�n:��1��I�4�:Ml�D$?��jſ$��g['���^�Ug�p/9U�b쭏�7n�+i<mFV���;=����JjM-Q�ɟ��Sk�K�\I�����k�z�CJ*�~zY�f�_A�����`���L��a��m>_�1_6���I�YB�y���q*X��O׿Wj���-?'�E+��cK	w�9�r6����Y&â�K��c0�b�^y���h���t%2��r�Ey��]?���q�� &h]��}���n�'F�7w*�f�&sZ.���L\�Q�Ҥ�'��f�RA�vw���MD~�����I�N�V2�� M���5K�i���[��;G!H6�n�����I�ko&Y�ff�!-Lڒ����'*w�z�t�B�b$U.%H�kK��]�8�*��f*뾸l��)�,�M���Y
�.#Ap\����~��΅9>i��oQ�h���F�+u$�i���T��8���o"�������V�t!8�s��:IP��E��X���
�2��5H�sg(�v^��Q#Ja�Ռ�6H�YDI��TE
ѷs�=(��l�,vl��H3��ig�Ԡ�9Sq�Ky�g�	��!?��މ1�b߿,Ro"�v.k��ǖ��n���C��(� ��f�ur��?�A�}l���I����(X¡��	�Y���������ʏ�W�`�R�EIb�m�*����9��|�U�6i���&qB��牨��Ѓ�;�q ��ט�����u`�ح�d�#쒼�]KcP����?��.>��i��R�	v���sN�|�)Y�1b�Ċ/����@�9�C��� *�����K��4����'v�A_֝v#X�_���c���{4��s�w*c�Ā�p�a�"\F�`?}6��G�b��x=����jU���Ū�������C����;hp�>���v`��+ 3�̘���-���H�S�f��t,r��ew܂~X�����u2c����۾.�I|W
�R��_����մ�b�5�b��p��q�$���+��ד�a����0v`��K�
.�Rep��;l&]�!?�7���g��
{F��ڼ�������yI�'��w�j��O��5��.ٯ$���N��T��.|Z�W��(������:0j��	��(Ɣ$�f�~���@8�p\��կ�[���D��lm�?��ŽȽ\��x�͒������G�4=/ 0tY��3����� !�I(�=��Ίj�)��J}N��K�y[�g�dަr�����ÿS�g��Jiq�tíJ{�����"_E�	�;w��L�A��j�F̔�K˫p%�V����\��ॸw�ݘ����s^.;��lq҇op���j�a�q.9#��-�Q���9����%��k����d���RG����
!pV���3R�$X����&��O��o���V�5��V[Z=$l��ۗa�g�0�`os�����B7��]�XhU��X��/W4������;�?���1`PH� �(lN)l�P�=�'(��e^��j�5D�a|�I��<��w�YH �D�"�7���|���Q��-�#���������}�F���ژ^����ѥ�`1�	��2r��2��ֱn��Ά��}rg�*X��P�dv��Z-�p�ȊsϪj���'��?e-�K)��A��,�9d�Y��G��LE�^v���ɂW�	�d�19J L}�uƧ�o��)��?9���g9c����|f֭�Q�[M��k��Ō��uYZE�Ӯ�̓��nT�ؠ���4�Q?�ʎM/����T���	}�{��������g8�$�֡v|n'�=1 �]D�v���j�]�u��8���*�0�u�X8�x�&�b���Πp!��d�q(GC�*���R�Qp�VP�s�Nk�8�/�aT�ꛕ/� �* -9x�]:J? �H�p��Ư�k����཮�`��3����j}��-�� �*�CJh�\�I�i<4�v�ۏ�����%Ne\�@R�u��ս��Q[�c��6���f���ϼ  _
k��g����� ����.l�?~;���[#�h���p�\�LX$[�\2� �K�i�� ����H*����l�H�\�}��ߕ%������q�f�Zei!!��	�g)#��-�R�?�&�C:B�0�y]�g��J�Q�K������CrEL�m>k�z��K��T�C^��Sy�0�����q��+b�}�BI��@��7/4 6M��
Izΐ	`:��$Sk�y���[�;G���o>!���c�����n����4�蟨ݽ���K�w�d��J��:��OH|�bt
.��l�]�y2�i���B=��_�%����H��J�&���[&���c'�#h����7��~0`��%Gܹ,�����M�ܧ'˂=,\=����N�*ۯc�����e��"�3
�ܨ&�WDR��1m{�ꏡH��gz�<����}1�8~�p��6\�֐�p?���!�וN�|�������&f������ t#G(}7��N|�������^���*�Q^���"7#��(��B+֪k�F9�-M����ߎ[����c@�+����|�D+���is+>�%B\�\d��ڷ��F#�grS��p�5w�D�Di�Υ� ��If�Sv x+ͨGD�1?΍�:��$ʘƹr��'�����Ӆ4�MT��$󮺏-&�Pvqm��S�MӜ
v_�/y��P%y.
0�����*��:�L=޽%Ey��6�3q�a�m�۷�1�d�V�
��E7��������KW��k3��Q�����y��(�^��R̲�1� _�-x���+u��d/	�t���}Hjђ����DR����hV�P�͗b��������쟖G(`B�+8$E(,�V�_�c$��,���9>by�m9\�c�t��\HS��Z
z��Unw�y���!�)��G��I��%�3�lP���m�9/4c�(	��qw��x�}T!q�t�>�s�� ה��,x��)��v>hjg�l�h*�~�+x�\��q����C*�m,�%�zqS��e3�@ժ�����}Ѣ�"�au�u�CA�ʻ�ö�������C�gD���FS�YWhq���ŧ�cӊm�;���D��&�I;��Z!|��1�HU��"�/٫���jr;s
�z�wo��I�u������ �G"�;^A�/D�=��m2���J��+�S�ݴ�����HH�o�HS";�����Ӓq�9�r��'����/9|rV�q��{�b5�ʥ���ʔŊI��D3m7���`Є}^��0?c ��uI��w>Gm�+��6���P6���w+��76���
����:��Cn��k�WC󼺺(D��>��kJic��ݾ\���#.�-�8@{g �|�j��k,;��"L�0@��qb���t�LF\|8���A�\�����H$e� ����f5i҉V�3kVRi}+u:�р�ƙ-�ebćz���QGG`�5�G��@M�AMK����)0
�34�IY2c��0����׿g=�M�>��_LH�ұ�7��ś���5c�6u���੝��?�v���[D'dg{��\��2`_A#��Gd�%���;)]���k��gۣG
�t�K� P�`ă�>ǡ�Q1�ϱ`������=�b$�@�J�%Wk ��0^->�h��*��0��yi�rɒ��M� |RP���AUr���mۥ$G��N���p$��0�oj*ͭ�o���=瞕/s� �~B��u��֖�'iT&���a��1G��jg�^E��g�N)'���-�ջ��%��`'+AT���"�{������.�
�X�����}Ǳ���V`c��3c&���*\�	£rA�KB����SY Jp�R�Q�5Mg���q֐�_���|���7���k�2����� ���$�xcb:wml� V�?�(��v3�(�ߧR�!?��UU����)�N��͘���o���0��rI�D��L�MJ|\�8&1�7���ae��QL��N|�+w�%E F�q�ȓ�1]�D��S�T+�Y��m)��X����dIG��G
Q9q�P�U	W<��Eh���2\�f�nP�����x����"���j�s�V�kO��Q���O�f�q�S�S[�`x��/����JKK?�Q�(ڞ�7�L��y+�U��CbOo���蓴QE�#���딧�'}�h>��D�)��sl�)��Ki�z�m^�#胐B����T��>��3���L�����g6qT@�
6��3hͧ�/��1�0�t��q�����*Đn���)�P�I���#���JvgMM}�1ⴣ
3�B���ȷ�(Ѡ�i�)��%�K��5C�Z"Vt�b��4��Mr{���(k�Ԫ�򊙺8��� ���q/��>��7}�����1y"%ы�ͼP�9�f�ت���
/�7��5:�Ƈ�W$5�@a<�n��֔Z�Bme���!I�S[5��G�#��ȡ��{,jb0\a�d�/t�&�@��[���|m�����<}��,�����)w�~Ȕ�#1�_/�Z�Ն����6Bp�H����G�K%/�;�NC�L�^�
V���!��?��.���^�=�5��
��Y�Ya�D����#n|�X�'y�F��\���d��M$6���̎�(C�Z��+��]qc���[��ċ���L���ws��j��-�W�L_��Nǚ�1'�0����㾬��I	�O�������H�j�� j�N{ۀ���EN9�v��ffP��m��NNtuV �>jp��}�Kf=�����,��Ab���!$�>��MV^i�PGN톟A�fX��=��%ݏ3c����������)��e���ckk�{��vS=i�d�l�+ga���ٝ��h����<~���� �ϝy|N��|���yO�_ax����ΫU�Uqm�MtԱ]���J�Э��q�x�B"�7�IK#���[�4���z��	\`	��>�g�D߅GVWW.���Q��������d�����"�!�{�˄�'G=U��gV�nJ������&ܲ�,;�8�gu��"W��fG�եnG�Jܗ;������M<�����@u1��C��w���g٭��1z��F����}�ґD"\t�O�Ni__�n��#�?�&���[-��`Z�iG?�0��^��RuUg+G�1��b��{/��1I�F��=iZ|��\oVH�U����o��]���^�s�=l'�ű6j�?�ͪ9cb���1n��6:�)��~��/�Uw��e��w7Z�q�5���kȂ-L-k,�,��a+~�3�w��<���Ҩ{H���e�?�Y�)d�e�;��X�����T�6&��Б����L:d�N�3w�%JDBHhh�~�<q0f�	��	����X����UP�������6�-h7ްO���jݚ�V/B���w�X��.R#�	�G��Ź��_�c3
!��	 ~@���M�%����uԆq5�
��� 0�WX=Y�4z�N����V؋*{/%��t��]y�)o�|Egq�rEJ=2�X����%�g9=��0w@��r=��^x���z�@��~4D�}�8AFzan{ɝ�Y7�N��#��+����}���IU��{��㹊�C�/�$��V��&�vk�-�ŧ��zm�G���b��:�=��}i��*�v�e��s��WI�_|��bP��Re�#�j5�6_�҂���s�-�ïOl����Od�Ҙ��s�r���̣��-�I����zc(������o�R�q�(��4Ɖ��K�t�b��Ô��ҳ��o�}����6�:gͫ �+�<��)�B��&���
7�*�O�N��|���������6��YƬx���OS:�w��O0���v���b��N�iT��\2]�*�s+��,w����A3��1%���9r�.F:'�R���9���L_Z�;BN(�'�P�J��ђ��c*�^!���2OYz�l�ȅa.	���1)��F��s����7_0E A��Wd�rBs �m�E�=��_>G����a����$�TCCL�� ��.#[��q㙫U���Ŝ�"�:����{�N��\�������c���I��q{5�1�Dz�Nk��+���\�E�L[Q���Ӏ
�G����W��Z�|���m�yy�cpd&c0�jEK#�� ��g"���I��$/&�l_5<��,��p>���GpF]OU)��v�#p� 4q=�	-|`�����9R�@��.ޣ*�zGI�d�%��B�cU	�c�ۿh�$v��shR,���\)�=TuD10-�J�tFB��^��!�J���i?-������w�-Ifg��$��l���w��o#Q����p}.��3P�b�c-�Wm�SeRKT�ǅ��>�*����?Jp������C�^��-4^9���S�i�����Aeh�n���\4�b�e�J����X�c�X*�O���/5E���~�c[��G` �:���j)����f��p��Z��ś����~7�I̥�2��m94�#��R`/�#V6b��7m�;�l�W��q��T�&�pR�ڵ�\�h��x���/.�E��T����� �*���;��F�Z�������6�"B�n�Y���6�3���rV�a7���.�`�DG�<�`�a����� @z�#́~d����ŲݥL�I�`ι����C<d�&�.&�z�~��#:7�n��������š6�3Ka�de����1yb��L�~�����c��{�I� 1(�U3�p~㧑����#�=��)�1"dआkۢ����Ԑ͋X�
���|��i�!��?#��\��Y�p|�x���R�����e(��<�J��[Ծ�N)1�d;/�����14�>�ci0��&���� ���u��3G���ߨ�2�e���9A���u�$�BVBq귓�(�E�P�v�Tȿ?�?Y�l>�H��2����[��X��fp,�Ǆ��O���(U�W81�����#�h�)�5��N�V�h޵6� [��4��q/Ə��K��E�hB-��,K��j���&�YI감i@�r��٥�d)�����|��f���$�8*�h�I��x��Fb����ZhDPd`f���A����!4G���O	 �"���an=$�V��iI�\��\q�@0�eq*��:|jW����0c
b���ܦ�A�����1[�l&�Ki���3Y��bVo����0�D:|����ZK�(��W���zN| 4�d����p
��yb�:o=I����MY$�NZb���q�~�%Ky��#���P37@$�t�a{�\�T�����o�i��dF"�њ��V����t燕�yx���9�$��O|2Y�~��=���u0�Ó"�Gs��p��G��W@z�����=�� �H)ac�z�;vϧ�vB�����)����jF%ǰ�DKӋ˖c��5`ԁu$�}�����^��Ƙ���c�T�w!^ύb�z}�nG�L��|��e����>ు#��ǩ��ܤB�/��sZ&s^���@��@���]�s��s2j�8��TQ�̖5<0��b@����J��m*�toBh�[��Ν��1����hgH���/�+�Qzޔ�D��y�|�Cҝ��lW;�I���j�?�Kj�.�5F ݰވOI��*4+�x��4Fw��������f\i���'�F)ix�/��t���V4�yM�	b��E��t��3F�u``����	t�Nz���[<󎾭-
6�x�5Ӯ�}M��XA�����P[8L�˨����z-5|D�sR:1�e9� ��]"�,q^�!]a��w�d�� �8�Y��1}FZ�X'S?Ig#���L ��T��&K�}�AS~����w�T�n`�TA�=ʆ�;��k�_�]?����%G'.*�@sH	��r���Ax�*+Q����2uX�T-�t�� �%3:��� u�1at��A�����)��c*耋�(G��I2�2��́��(<�@�e�{n�nxL�	�%�#M�5*v��z(r8Qѵ�Ni{j��a�ٮ*��l��,�_�3*̿�v#Z�	��N�)T֮1�Ǐ>�����.x���r�p!�N��v#�`>�.���_�޳���ba��2Ċ�������6��90�KC�Lg�w_}U�I(v�#!��� �u��ʏ�U��b���%��n�/�攉�!7�Us��P5���W=�6j�]~�+�^{�~R�x�Q���J!H�1Q>d��pr6W$�5��w���������:Ԁ��bV��O�6����3��U[��]�����W�c�'{���K!� ⳔD!��u�ȃ��l�X��l�����>c좞0kjJ��� A#������v,�㝤̟�kNpB��SK+u8�@E���$������B��h5����EmZ���oą���/O��_��~oBН8�5�1�'[��g�L�J��uՆ�oa��6S�gm�\��=��VT�I��A�\��;K.q�e� @��}�f�i�L�@���K�7	c'��C2�bE���ݕo�qd�X����ȗ��5G�#���w�ͬ�[��T�;����Cq�w�~��*�FRZϔ.c�N��r��ܸ�g?l�Z�B���}�D�uk#є:����Q�!À�֞3��ձ�g#�v�z�xE`A�Y÷���7`��88�Q$l�Ko��Rt�ќ�l��֒���4��<ݼZ�C�6��F�o�n�;�ȿHk�-y�'���}��?q���q���5�+�B2�y�����	X��.[W��-���0d�����T��>��i�VG�ꁼ��w?��;�Sq�~M��V���"�2BF���y��Ϋa���b�_<����?�����Հψ����~6�)#��i��o�qQ��D�$���D
b��~ח��<���/�ϼ�߀ _�\V+=r�fd^��y�a�x�� �K����"��`ȇ�a���.��2��n�����22K^P�Tg9�1G���x��қ8�q[43Vʲ�s��AK�=�X�M�~�M�]���Tzs�g܆х�H����딈9�qz�?ٵ�*d���/��>�V�u�t$z�^�A��=�p�r�)�1�*�p3��ǎT'�8����dUQ����0���k��t�	��@2n�=���+ddbkB�#U��b�p�3��� ��>���P6k\�2՗��������=|�QÔ%~�.���Y����U����Ћ�b-���'z�P>����$�8�uK֋����GK��^�~�,^Lx��a�O�̀��˔a���7O-ۜ���&���p��ܹ�*vR��$�N�,)#���e�WH����O5�WTר�4Hc3"�A�q�|�
��x�;�m�����=�"?]��S�����	p�N��h��CX@z�$`����x/���e5�gV�f���/�f`gH��s=�q�O�f7��45�ѥ,uᬖ��քn�+�9�yY�/���=�.Ż8lK=�#�x1���~l��/�/:��[��E�(��Z����O7�,��l�=�������7�����x���l�������
��+��8���%0��a�~����1��T��^��q�H�z����P;R��_#� 
"U85��Hmz�"i����N�z,;F�B�$��P�Tl��� ��t�DQ�^S��5BL�Gc�׻7�X�C�&�3zw�_�!�l�z�q�:YBO��_j���x��L���:�}$�u���h
Yf�n�ϔ|.�u��)��H�(�D:��~AEl���Y��a�٠k�|(���Z�]/�q������#Eu������i�z��D�H�e�)�]�n���\E�>�;����IӒ��{ ��h`>�L���KEݱ�ְ�xeg�$o��~����vG�
"�t�=�y�Q���A�t� �
UWFF�O&���<p֮��՝���a"�.!�+[��i�Χ�N�]s�6�l�{��F�%χ�^�}��2%��|��t��iYg`I��c��cS,�?��%s�E���p!��g1 ��&h���{	B|�0V��KTk?�'����y�x�r�8��(��t��::�"�kr�r����=����ފ@�=�@H;���Z��a�����/>%>H�}�"ƞsA��U�B�㞷B�7�����>��۠_�z�"\.���N�C.��P��ڙK`���eՊao�ޗL#��*�QZA���f჋,�������jD�g����,�l�m �#`�d�G̐�v�ju���zsP�++���(����vZ���Zo�2�v������lE[�J�RP!�=C���<�dd�w�>T��G.��_y9*/'��Q�����$��n����N שFmr(C�],\߳��e�l�tB�^�2	$�;h���T �Վ��;\т��;j��#k}A�a�d�67�-q����^F���&Z��V�� #I���ڈ�bR�骶s:k���LW}������H��-t�&e�D��:�A\�H�2��hh6�$��a��p/��_i!$�G,Z�v�پ�n��8F���o]�T��G��0�����:�b�m��1�3��/�V�=աq���.E�a9\
Fn2�]���O^�$��P>�<%`;�.�)��a�ܑ�	U*D~�\��hg�I��
& y�YF���;�[��/�1\(1ʫZ��`�Q�;Àg�8�[��z���[���g�<|o-�B ���@����&-C�!��fҶ���0��O� ҥ��á�-���6�%�P���n�K&����󱧳i�srb$�l�8oޏ�:��{!W�O�Ԗ��&rnt��yK�i4�S�n��]���Wf���C�̈t�-x�~;1��4v��v1R�t�|��Xw[Ud����+7hzk�����T܅�QE����腅��+�H��&���٭2ܪ��ܛ#�Y��i9͢��;��^F�蜷��:�W��s�ۆ�a�5$����J�Q}o��`m$&h�t�M#�Et���;5'���s'Pe�&F���&@ BT��^�H���~@�L����E~��������w}<�-z�	���ݼf��CE�><�v%�6gsz&����c�+���|M���LS�Z����,:+(Yo��y����"��e/�,�N'����/C��ĩ����8߶�N �+^�-V?F�6l
K��Z����|�ӟ���y&������tXz2���jȺ]�t8x��W��r!�-q:��yu3զ�I�U�D>��1���Θ�x�=]�Gq!_!��ܸ��k�Ώ�e���������#�'(��������=e�>�ئ���N��sM���Fڹg�Hs��Ȍ��Ů�@�z/��Z��WĭĨ]c$赙��yd���d�.B���-h��jT��3�L^����O�M���G���VhlZ�
2���p�O{3w�A^�h@<��T��Qw��c�?��&�ـ��q� 
z[��<�C�����>x��¶�<��R
Z�V�E�}�C>o-E
�\y�Kh���.Apz��M�����r;�r��!�uNihBI���LI���zEj��nŬ�9(��[�u�Qw�F�I�����?�=e�?�Hㄌ|Za��H�wi������FP��b�4�ҬX恉&o�n,�PN�`���I*��_	���Ht�����L�4��jl�����I�&F����[eӿ�
�q���a�:,3O�R���|K����s`�8�3lZ�*o��g|dI��Zrƃ���f�n�{���n���P|���6̐[�+_���L�ȵn���."�� �jx��%起�\��0�W�1xa{��5
��̇������ѽ&������|1y�0����,�#��1:UM�[֍�7��
�5�����H_`����*�,�N.����rG4�b�qJ_T}��.JL c<Q扠�ċi�Y�v��λ�7���KU����t��]��*��{j@ٰV����y<Q8
�0�oi�)T��ݎ*|���[�[��in;�L_W��o�%�xRŒ�b��G��ff�lS�4Ic,����r�Z�~몢.�L���xG�A�WdK���Ul��O����
_��^�y�1O�-�5b��3�^a�-u��j�qH��:HϽ�f�+�$�H�2̰��x�Pܹ$6���s,�D���G��Qk$YkT��/w�����*(9�xY �������<�4����^�������$���J�����%�#���=���mQ^4��;��Y�x����
l�b�ּ,Dj�f�u/N��-�<���Yϧ���Y�}���NQĀ1Ұ��/V�zѿ�6,��������,O5��|4���G�� �n�����xrc�-3�ޭ���2�`.�jD�{D�Z�XT	��1 �M���@iI/g��\.ۙ��NE&����=�AJ'�- �����l��e*��~mx�a�����z�{kY�G��&��6/��݅�i��Ϯ�vD���o��_��"n+2���4������l!�����V'N`#ƒz��겴>�"��k���$<;�D�h�����ꛏ4y6Q/���/e��4>5Ph�������9�Ul��S�Y�d"�I�]sDgڼ#;(�l_��k���DR�ʋ6���{J��|��O�"�N6��v%�p3s�$������1�(��T^��A�@v�sఘ޺{�o&�먴8�4�`nB{a�H���v&��)�~4\�rmV�����q2�{�N	(AIpjM�/��mւ4�GZ�\灹	 �~��Tв
;4RO�8������}�Xb�b[�NmVt\��=�)��~"�9 /��g��kk�bw����\�����c~m�������@�v��p'"+�D�F��< 2�)�JZ�q�&L���2}�nL7m��Ȑ���E�_n�q����/Y�d�D�iJ�\�0~��m�̍ŕSt)�k�C��������⏘J91�����A���'S�8�~"���2��=��G��-}}�해k������!�+��P~���З�y�Տ�����i�@�q�x�^��W�zN����*��Z
m��(��-�8�5��;`Z.?���(���Q%����V@�z��y�ʗ=v��S&�I����S�i��� V��!�d?z�������qt,�16h��g-\~�������0n�nQ�q"��g��0<d�M�/�9ffo����_���֓5�]�<�~��]q�F�8XFEM�70��UD����Іyܭ�{)�P��������M��w�O��q5BA?���{���z�����1p��aؒ�G�f4��-! �'E���t1C��ͨI������F>�����+���d��Y�wΒ�e��$���rP�_S��`J��@��//���*A�������Yo���4;g:o��]�foJ��y4�����)��#d$�@��uO�ً��� ��)�'�8)�U�e����*T�/����=�Z�`�!��c�o��
���_9�*���]�g�������X���~�㛾�+�@�ך[����Xit B�#}���q\��)6��6LC�$~~p�jͮe�d���U���P_(V���$��]�7zTQ^����
��C�ݗ�4�팆�:��pJ�l��G��[ ��̈́�����a·š����
&�-G�`&���x8�lY��.8��2d�q�i8�����B	�y@�,�l��?JM�M�|����[���Ὢ(�s|/��"��	"/{O�1~[�pGea����_3��x[�0}�i�NiA��M�S !��\����1�Hѭ��o�OB�a�^�I^���f\ݶ��D�T4$��Z�V�MM�r�"�:C�J���+�o����$���v��鮞{����������ƫ��$Na(Q�J[γޗ[�؂��33�9��-�{���KP��쥔! A&$O�Q��ޔ����¶����)�qs�n�@�X0$�>.���râ!f-�� ����LfP���-����X�8��"���4�me p)�k$~ߋ,3�`��Z��z0P���� 8i���0��:F�K_����)��V�qt�Ec!8]�;��X�\� �-�{��H�"��7�ú��g~w�q�QK�UK�m��\��|*ˍ,�p�b8���ʁ\�
u�k2|���/� �)R�U����YM�P�ږ�!�:r(2��m/��"%�?���oj^����hC��E2p��{��EtgI݀����~sq��C�o��u�n�B���q��i��babGԔ�\��:x�[�?�|��'W�yp~3R�Pq�M_J�!Iͪ�T�.ެ5�X�ީ�1+�`-WL5�h���?�]�Dj`������Hsvb'յ�4���@-sw���S�i��:\u��\%�h1j�D5�I�XZ�y<C�*%���Eծ_5 
9�򂕃$�N�#��)<~ �yj�_�����n�>�R	5�y)��R:��"rd�!���U��Q��i���X�H����^Ҕ�����	1ь��\^S�&uԡ���m�W+%��1���f�)���!��ԫeb�=�}�ܲ?N�5��?�n��h
�IYjxJ���\�L�I�/�O�S[fc�M�M�w|�j���?^�^@�����7��8nC׈��d�T6��E@+)LO���n)w6E�{�o�y��K��.40Dg�P=W�%p<�I+8�XTD8xaY
�_:�'~��|$��g��ۑ^� �)���MCMny��똃��
�B�Uǵ`'�+����<l�].�܏��t@*~��K��h��	n9r�4��	�p-��W���/�i!�$L?�h��Y�����3f(�5>Nr��,&	�1�!�.�:#�G-2(�.����e#v9 �f�S�"�)>XY�ar��9�o~�Ǟ�J�����u|��EV�w��u����Bs�'�4�~���uI�c.2 O�V���7��[��y�&T�ʹ���}�$ɌǦ^����?@�FcW@�^�Y�����Fd���c�(�H-Ɖ��I�MŦ�!�t8���%�72��T���r�A�%���C��ļ[�I���+9��$:��S��+=�֐������K��� �ȝ�4�+�F�4�!M�$�Eybľa�wg���y�8r7����h�Hę0��o#t�H�e�;��g�^ ݜ.�I�FSF��ZYS�s���&?�ZjF�	�����Œ�F�齌�J�+�ʀ|K��#4�rcو�e��Q�(����mze���|��� ��Tǘ~!�O��3�Lh-*��q�1�j�A�|�SG�4?�ke�i߂s5~B�7�����!VVB|ݞi%���o"D���ђ���wA��0cb�#���G�0~�A6��C�o�
v�0�z����|���K�k�_Db==_ˊg�����]D_���t!�L��oD
gH�ߊrY�2���Q�=`A���A��E��P?��%��Ҝ��O��)�R$��-��T��1��g_?5;�����D�/7|Ѣ�[�]{}�7��Kj�Й�#ť����̫��A����{��eXs6��K8���rKn�TT�ِ�<ZG�0��oe��c��WN�
H7�S �/�!Jb�p�LZ^�3,�
��8O��z��zi���E?����VPc�&��{착G�]�O=)KE
'�ee���}՟��5��Ā�f�A��H�sY�#�i*�6?�Cr�� ���[ܠ��	U�����b</[�j�O�ʡ\���s��mR�o˷~Cn��RH���rY��V���ʿ�}��:�=��S�?b��"�iX���G��j?/�s�� ʆ�G�]�Ǵ��n���w�w'@R��\~�Fi�ީ�b:1.{!�I���<�C<ɫ�}<�7eݚ7�c\�#��2,����g�J�ݥ3vӠ�πG�kw����|��)�����14j��>y�s?Y�8���wG� z��r���x�OI�*�|"���Gm�C.��%~㳃*=ء)����GA�D���N�?��*p!brz['a8�P�4�����{�6��c��IM)�h�����x�7��w����B�
t�G��5<���W=H�kϥ��8844�u#$	�DTM�tD��f���^��!V5H����#����c�]�u�|��=�U���h��e��|g�rPͽQ��Z·g�cܾ$P�M�-F����6�&-=��c�{p��:j��'��20WaC��,|�/����r#��j�6č���hir#'"��U����9�/���A*�(����m^Eo�s��-�7�/ٗ0����YB�����W�:��r�����5ĕW6a��O�-2-Q����,m�iU	��u�*��:k��q�P���ψAP;���9&�{Z��?B�c��jxC��H�*��/i)D��|�<��' |��2w
f���O�1uVK�H�wt�3�d|f2a�݋����Bqt�k���qڴc��T�Y�p�����8�j�@Ј�ɤωx?���_@��JJ���_��c���'��ðy���&��@�/��Q4����^^}�p�t��1��o��w��I�^gF�|R��#	���yܶ�ף�3r2�g%n����{M�4:
]�ޱK^�<�Wq˖��k
�`]�|������<�D�{,�{|�����^Բ�}��ca�2Т�AL��3c�x���F�p��f�͉�C�#��s ��X�p��a���Y��U��.ȽV�VG����=�7%#f�L����`�Hk�Yʏ��[�h9�lԔ�|���s�I,��y+R�̵����L�gA��4���sA��)t�Ev@��ċ���8��oA�@����;h=�a�\�6��|Gu<��;h�Z�L�.��+�C�z��4k,��ςS����e���	!d�m�����kCJ����e��g(�Qt�u��y+��W{겘i��zhS B�t�7��
]�+���ͩ��4�H�/��r�.��-�w���k=?o��}�Z���냠	�a-ʿ����83�9�j)UP��A��Be�n�����v���I��6��Ӕ���r��d
��$"B#����2!<�
�%V�� �p�>�PM�������,1t�tJq������o�\�#ڒ��������Db{��^b}a6�ws�z@?6`�F��C�h�C1����`�;j]���������0ܒ����Rώ�2O�>Md�Z%�˞HwZ(Bȯn'����B��bV�N]��Y�:NW5Xw�'�n���@#�u~Y��gj�/n�ڝx+�Kz���f]��Q��hي�5�yh�y����)�/���]}ft�XR�bAy��(�j��-�J���-�g6�a��#Ȃǻ$[�v3�����BB\%d)s�f?����s�sK�_w��U�x����\z�㚺��e����0j֧� >���tW����i���5b���>�'�AG`����x�N��O26�[6e?��!�L\�E]���'����I�qug���x���*�+�ܺ���-��*�Á����q�Tb�Ђt����/.����u���4/>ϭn���XӸ��c�h)c��~�2�1�J��˧�L�M�Ȥ� Ok�E��=�����&�5o�pR%3��`�8�_��氰Ǟf	�֒�	�t��m��i5�q[��G��6�b��`v�֩G�0ԘI=`���
�q'�)Q�	|s~U�\��䔎��.Y������0r�]�F�8JP��s��$��H��V�Θ��
(��� ������W�?�.ٕKT���L��7rw�#p�#���5m��|�UDv��+C����%�D��8s�7��g�L&�+���4��Z���(���\A�Wa�Ws$�C���n�/���ߚUBU.	� q5��`���ski��,��K��N� +�x��0U�vb77�`���*�Vo�t=�(t��7��7�� "�N�Y-�(�L��ԉ^��9gw�C[}��#�����&y�;A����d�fr��<��/H�~�'�Q����RMX�m��	��6hJƦ��Ǘm/&�ZHB�o+G����n
 6��P0"4oyw���'��o/�3������z>j������Q�����*p~;���Uz|l�"탼�>4�`�-��3hd�<YTZ��|%pi��x�I�+�b�3���\���g-��ȅ��#|</���o�<ʥ�Ҧy-yG����NvC}��5�ۆV�߇���|��[b��iV���.��*�A���V9%��)fz�#E���U�����k�0��Mhl��� h���ɹ|�q|�>:|�ٙ������9~L�'�����Ly��_H������w���4Wѭ�����>�5B:
��i��:��׵�(���z�yحz�܍E������ �I�����I�'b��rf��v�W%����	�d�ԋ��b���O��	>&�T#T��
�s�ٶ��}�Qw��JL�N$=�J��5,������R�m�=��F������NiL+�J�wJo��h���m�����`�e�qn��!����9�[/��r��h�υ�=��=	T����@�� ���H*��V+�Y\���K�X��*�8��7�W#^�� 4�V���_��j��r\Gmǆ\�����J�kO�ʲ34��rb4�X��'�Sx��A��k�l[�eX������:�㵁,�L OY*�4�_����_d0f��JIQX���8��R=5A7tgtى̆��W������(���>�D�VQ��r���N �;�ܖ�����r���v�ӷɇ�M��_yCm���]�&٥��a��$�4���;��BA��D�e<vkF�E `�
�,��k�tW�����d�#�4��z���^��9/OR��Ê\ͪ_& ��� ^���U	�)u����|�V-k�i�]��i��4j�L����R�e2|�v��[\���t����7򒘟Wn��3�^���[�~a�W�O9���Lk��@Pc�rF%��hYE��}n\���5�^�Ü�g�H!1��#�I���'��B���XI�o��~ޔ ?|��Qs1��`!h�\�i���y�(A���s�Fռd�5���&�mT|S�5�ImY����X�Y1���c8(�	5�1.����V��	���n����,ا��T�y�j�����<^�@���l����2Wiy�
j�D����`Ҩ2��M�Rϐ#	A9'�%It
�l�P�NF��7-��>1+�8���? zƠD���fxe\��b�Fxsc:҅��:��gp��'���w,f�$���^�����g��=��4"�a.�?��;Z^��x�v,�"�m����<lV'����`�A�'P�KA�i���T��0��[H�J� ����11us�����o�Rɉb��"C
��(��j���wt���`�nw|v�6�[�]�oez	��i򫅗�c���ǫ ���}�_a5�+��u��*m�C�I�:e��:�(�1(��_�	���8�������3?�w�^v��(�#H�6�H�6q:_\����å�����a
��t��d��TEM�"�!v"�~��8�ҬY�gC(�߽#���H�R���g��+���Ҭ�Ev���;�n����2_&�	7��.+7��@E1�tsR���,��QAj�n�����7*��D;<[����`W���;R��6�E�fiDB�nkXFz�.�$�-��&�lyt� ���D���ߓͲl ��𦭖�$jF�5l���Sފc��[��6��Ŀ��v���Ɠ���-"���ݨ��iԷ�՗̗����Dz���%�3��	��$�Oٌ�0}�f��p�Ʈ�'���tԌ:�7Pw@/�:*��m,�.�eä@�:(ͣnv����X��|�����Xڴ��|Z'gf��S�U6��*����C��B�����ڎ�PZ��Cs�U`��w�`q�m�u�Ld����W" M.���ԉ����,�+��p�/S�wB�����z}7�?օZ������ �Vx�Ꙥ��h��q�U2�wQ����=Ҟ�D!J赋-��װ���Sk������=]S�k�I�D�����ܾ,C�\�T�p��"��z�W���"s�u�?�$�0�Wa�j-N^����C�t����Y��k
�[tz�3�s�%�2a���P����+�J�K�{J��x-���Fe9x�p��|���(Fl�2w��D<*���dm�U8q"珞�X��X=��.��y�}�QN�s,�����2n�@2ڽ���� �9_#EI�i��-��u�������r���s��e�*�-B��'���"d|�{�A�R�Xd)�A����Rڹ=i��im�Xژ#8ѷ��l����G��i}j�c���6�����S�#�d?��H�,��j���*��P��JjU��bq?�_'Q�̇�<4���bp��͋c]����\��'�3:֤W˰�?CN����FY:pp՗��l���btj��:&f%W��[5�h�HE�)0��t��vY`p�.,x���4�7�[�W�k\��?�갣�2�5��z�m�k�|� #��/�a���O��GWH�K��0�Iϙ�adzy�Ph�Ny��z��Fj����6�"A���-�"U���ѵyVFx�{cc?:���4��_��G��S�E0���Y����!�&���1!�7񽷁A��������������
���𭜵|@���Z]������_8���[��Ej6�q�,�V�5A�(y�g4Η�(t�D�Sf���+\Si����дD����1�r����L�[v��$�\A�}:��n�vUA񲕒U�ݝ5�ǔi8B�s���uj������Vם�����c�`�Y`&�;�K���}��Ĝ0Y�"��#+����Z�W�>MW}��߲)5oI�z.������*<�SV��Fn>�A�Zl�y�^�Y7�����#s^~�kw�� ��}����A�9,|8k�ˍ��D��V������;Ɨ�E�a�w��b*"��Hݩ�pQ�����d_�(�!ڛ��7a��F]8�ka��F���9*ʠ�&E�ٕzd�7L��ɩr�X��F� >7�͖��� �=ň���Kh���l/��:_���� ��b�"��ȹ��M����l��ܣ�p�UQ퓨n����,钑~�1R�M�8��!�ȓ���%rv�&DSZ���E��.Ֆ�{G@�����mi�4i�P��.��|�hn�,�U���b�Y�s���rU�K�#�+$ۻ9ߧ�4T+��┵��a؁p�'3��$,Z���q���z� �OT؝ ֖vfe�7� q�˘��9�t�6򴵈�7����"A��Z_}�TAfZ�l�Ҏ��oKn�2p��&�hws�,�8q�Fk��0��d+�;����8w�o"�P3�J3�1����6A�Ǌdǝo=ca��[���5��n-hh�?�2�A��e�=a��'c��ɠ�����NTna�o
(6Z�`S�Q��PF�:�3����N5��s�҉#s]���?�q,6�U�@w@������mc����	�q�V?���Q�r��F�PN��_0���N�sv:����?�]�!�*z~R�p�SI묱�1�	�	̭,�Ԥ�kT�92���ʙ#�D��S�w���3>��8.T_n�q,O|B�Y�e-7:(��Ϡ���
�����p��HE+�9�mډء�&��{Rőa/�Iɟ<� �f{��"㭢B��[��*H#����?R"�4��0����x�0R Bl�62��<~����K�H`#Ns>����X��˟{�7�|����pѰ�g
/��$tK��i�v�<�X|Ş\S������.�'7��G���:m8xNA`��n�����2�������7���M$�j�o����c��𘃅��C:y�:�ϩLp�d�7+�G8M�*��46w<�y��dџn��|^��%N�:RcQQ�����h�����8�)J�
�cMv���l���yI�b���
��A`���Edjj	��g���v�w��D��آ�v�<A׭|�N2����+���+�	��g̏��:je���f�|�%Z�\�M�u?�j�ҡ/ߊ����5z�U�Z`��G3�U��w~
�4kRk�z����3d6�"�l�BF�����`��Q{�u����	�NH�3>�Ci�H˅_r�OR�4R���5�%�[��Z�Ba����C��YX�HC8��x�"�ؚ6<��"~��hk���G�����	B�7���/kt
�i{ �v~��4��[YV�� U|(�1��[�VSS=$/���ᖥ����J^XU��B�2@�X�4�8[�p!;fI5=�1~�|�_?Yc/E��kBf��gf�����A�S`��/!{z�u�B(>�^#d���=��%�������@Tb^$ ���\�$^;2��������,(x�P��:�6�>A�ba�V%���i�D�� #:���
1$��B�,���)z�l�˰�o	$	-;��V�cN�0�{FA�m'���]C�9[�Mk��c�,�TE�3�S�U.v`Ij��	؅[2���aSB똶ױ� �E/^5 �� |�tG�~��.H�����A>n�+/#��}a�6�{=&�*��t̴�c�|5o=J���ٶ�|W������};�-C�t���/�$F&Xx�Op���_[CN���:�Qr��єy�R����xR3�n�;���g����/˓�EC��ףM1ۄ��!곡8�	�j�IIx%�;��Fߪ�_�@d�����	�
�A��Z���`���(���F8�ǿL�sL���[f�r��v���.0?In����ﰢ�!�_wU�&��Ɗ�jAq��:�&�P��cg(@���SZ���H*oDOl� ���?��.�����HO�g��k'g�T�,v�\|#��F����TQ��2:�2�N
E9J�~P#�'�(0 ����K{($�r��s�s{��g��������p68�&���~���D���!4�dy�+"H�vG7�:Z���6����f�)ۮ=�pe�k�f����{9�����Cn�����-�R]�7�Z����ĕ�rq.Ԛ ��@�v�|��2Xo�/Ŷ���{?N��&����F�%������\�.�L�]�˰��n�[��`S�&��jM�;�	�	צ�?�)�G�2�1�2+7!B��/�-7�-6�&l	�/����ת�T�rFg8�h\-��ܫ1�_�1'4M�S�Տn�q�t>���p����"D�-��18��n<����i,Q|]����mD�ԾT�$�6�K�|N�>s{H�����O����gP2��o�0	u��A �8*�xOUخ:�)43�t�e���>�
���UyG�Y'�����Z�(%�M�]t�Jh���4����Ĕ����YcA� }��T��=
��l/1wb_�JH;� iS����46@�x�i����k��s���ҭajW\~��O����*M�^W<���B%�P�\�H�E�U������x�X��u�3=�to{<1yUmA��&i{
��k����V
�Fh��=��%{���l��8<'d�Cu�Ud���R�Ҵ���;�Xnv�k��[tz������)bJ|I��e�����$�%5�`=H�ӝغ�9e�f5~�� �fk.\�W�Z��? bg��?�\����`,�C+�2F$�nPF	�����p;+yv��Nʥ���@#e�R���R��!@�vH2.�޺��+B�/Ab���(���N*g�������9�Q}/1��V� �Ap7`>�;r�#�n�@����V3,��s�x��U�E}c��2&q6��u�u�cz�b(h)�9o/��a�C r	\���
}�̶�9N��hC��ƿ�6�hy�5-YQT!�a^Wg��s��;ꣿ�����N��z�T�,���.�\���y�s5~�v�h_�	��GVgX6����`�`���֢�F�������p��,\�Wl�K�YD��h1�$~⣆�"y�ECs1F����8ش��������"�����0�m�);�Q}��?�CZ���4
{�z���n�s�!ʔ�(f�� �ʓ��	[n�5�$H���6�@�a�kU���{>s�N�����V(p�}���<s���f��_��E�JR~m�ZTl�{�u�_��$����q���еM�s��(2G���7YV�:��Αd/)�Nk_V~v��e���o�/+/I6g�UF��J������������{���k�*(N�����d�w�M�g�kպF���ώp��v@M�iM�UDoL'�H�B����ޚmdQ~�\r6����!�S�`�C���)޽�a��鵕�NZ�
e�H�Fɢ��j矐�ք-���{/�����؆#�]������s(��^��u?��~�,�Z�ߡE=Ь83�4�_��b�����"�d�Wk�]�.
9���W��Y��lu��B���8�Z����*C����e@�L7���j�y�ɞ���?�s�'nd��z����i�UKv �ޗ6S���I[�sAI�Tߜ�}NRu�uo2Cc�Sw�D�ENq[ܘ��ۓ��͓�&eY�ɰ*o�E;��[)��t=v9��	+�eX.ox�*��Ĥ�h�_�o�n�H�R�$/D��o�c���x�viC��,�n��e���
y�2����/Z�G«���Ħ,��mr)0��c�CYV[��(�Li9_����v�.����<���u7d��S��P��D5�c2QZx\��&���	T����~�#1I�M��ѩ�\�A"w�=����X)j �S��,���ue�Ԫ�%����o ^P�&�R��=��8��,�߻~��<@[�zL�KeR^�z���*���q��攰K�2I~����&�. �Qs��X\\i�WX���P^��%�!�ƶ�G����Ń�Fj�:Gc�ʄ�a�E�ן�Y�� ��2t�~ 5����y�$�	���0�;�s�ZW�|y�[�a�����d^aC��V��~z	49�&�_
�!���~,�����k.>vD/���p:�.~�$��^&᮱�˕����ϲ�,�D�>�I���{��V�H���2�� ��z{�' ���Cͱ�g�v�|Y�������;�$j�N�ǲ��^j�h�1T�>���Q����4M�^�	;��6J��7�t���(_%>��`��<>��l����ӛh+	.Z:�d�q�X�bίig0s����VFX�J���5���[���/���������d��þ������) 1b��]\�������FJ_/(�W�IB��~��Fn�������q�����d�8]z�
}9P���I���g�i�%cN��?]�N_9^��ʛy�(�c��P�F��Y�Wq*�p��Ԣ��z�9��[J�&#׷K���w1J����a��V��Td��8���}պ0Z+a1�-_/)�7h���j�$�������ᨭ)�gEJ$�����3�z�TM�Xz�vYοB�`����h|5�7�:�aETC摅��a��J����hȽ�vv?�ۼ���A:ݐ?#�Z��n��o|K�)�.��+��su���!�١���j�B���`CP��1	��x�ŵ��.�o���|��:&��3>`�Me��N���^<&�ȡ���f�W|ն>�/�EG��݂=5�ϞS:�0-�_~�dVT�|�Ns��ZG0�қ��R�չ#q����`�����. ��N�A���e7�T��yB^\�h=w�Y�#x��˭taH�.HUU.��9���������Op��#�PM�g2���^��	m�����W����8��&�a�".��#?q3�k�ʐq��?-�8�Í"kLs/��8���B������x(�AAؿwyfs�Ӭ�ح�=>>��~]m ��**���>VF��-�5�
Zc��c{
�P�P�"�̨�Y�Yv�Сmm���L��Gy�f��uxc����$T�"�%���e����:��ޥ1~��]�I�A����S�w��迃��O�KM΃g,DqNr��9Ȥ�|��m��i���಩5�P���(ö��*���w��Za�Au�4��eq�3D	������ξ���{@����&����ԨE�\����DrU0���5���g�T�L��c����q~/�h���y9Q�Y���+(��n�5)1~g�<�}�;7��~�3��ua$� �Y��9��� �^��?m}��M
F!Og�$�l��姰��{��OU5i4�S`0��ᾼ!�V@S�k�M�y�H��+�kOq7eD(G����X�ť4���$!����eʏOLJy�8�g�uu6�a������z��}O����(
n\L��@ka��j�F�����[j�yI���c���q�VC�ub��g��H���	I�K"+Z�a�-Z}�<��N;�l������m���(b�InNohD��EN����_����-�|	N1�2
��Ն(��<�{#�G��)�kR�Aܿ��D;��Ɖ��־n���ch������.���|K.�>s~:����W.�?esGbc�T�����=c�����O,5�a3��/N�� �'�d�^�㳗<6"5Vp�"����Dˑ
O����Y��<�ɫ�9q���$2�1
�B��f��F��� �X�Ȗ���}��z �� �N*k�(��!�j�x�L�����'�`;,g���Mkl�jjT��Z�E��	�7)�q�Jx#�+�N@�6 ��$_��;�A��^lQ6�%�2��*�m�U��Ck�\�8x�� ;�iN��UK��O��+.�Χ��)%Z�ne��hW�J�!j5�=:M�LsmkFE>����s��6?���G�ӈ�i�9�������up�q�k����c�W��Y�(�қ��}I���]���S��.�_pC=����n�!gk*Oi-����㷖�����T1T��xV��"�I��m�V��!���,!�Y[\ ��OY�7�^`��<�0P��X�ie�_k�S��(7�E�|��+$��q�����/���Eem`KxƢ���.�3"��^ͱ����p=��:�6������K�h��e-B{K�*�b�8S�Q�������@��Dj���{��X��7����5e-t���fh�X��K��kFk� ��IA�ܰ�v�:�x���zڟ�q�'�u�o��Ƈ�rHv���O�1ᛑ4���B���*`���;vdeDm�+�N��3��HJ<�ܚ�{c0�[w��Uכ�{����!� ͠n{P_��K}s Yf߯?�5���=���=�09W��vg%B��xc�)�ձ�9�C�}�*��S#�#m�7���x�һ�aL�n�ҽPӒ� k��R�rC70r�	"�
��ڵՇ'�;���?'be4�\� 2�7�/�x.0�yz�=g���~�W��(U��1�(�ڪ�w8("J����4}�z��ַ@0Q�AfLT�pB(���B%�q��S24�^�R�"��ƙ��r` �%�۝мNt�#[��N�z���4wQ��pU�Q��w�C��S2��r�e*wy�(Mģ���պ�@6D����23���	G���	�5J�͜��h�>��sS.�5�3�(��e|)z����t���%��&Q�� �W1^��l��hwʬ���^�Iry�Kw�c����\ͥu�%��p"ŃË�)羶i���:��3)$�_��ĐN!@T"O����ez���挧�-�!�"������b�s%!�sʦ3� n��l}�ڣ�;��_�;�tL���6����X>�%�VM��]X޳�R\{��?B��7EK���%.�:
�`iOo�Vp^	@�w8�t�\fMu���ϧ�j�t�Ĩ�����@LS��E�U�x��ᒹ�v�F�y�L������]f���m5t�
�{�����N���� ��>��71��w�#�V�:ݗF�:�+�ﻌg�C��!���3q�3VX3aN���:IP[+�����<;�a��V���m�oe�!����+in桓����u��㇫�V��
������"`;?�+!$Е��2����0_^�7!��	�x��Y�{2� �XW�U��d�����.d4�ꠃ���|���:<����1��C�����L>���݈=g\Iey��z�,��<���9X���IA��"�xk�A�l=5�����k�	�r�
0�I���ka��TZ����bFYs��B�j�A�����Y0g΢����l��z��ڦ�}���u�D��W����1[R�	j�iD!9��[�`�o�9���X]dr���P��'3`a�hi�>>�1� �\8
�/�$�9���WqV��&!E.m�e��U��6�Op-��Y^ēc���X���r��Q����b$�����?3o��M��{2P� |�rN��i�����b8//5m��w�C��L��^��;߃�%&}�&<?#�7e+�m���� ��t#����i~E���jM�ug���$_1�5���o�]��<�ʻKN_N�w�����4-A.��{�o�N�<*�׃Vj��'J��y�>c�C	J���-�����- s���Mdq��Z����ie8
<��tC��g1+�E�x����Nԅ|z�+yS�/�a	��ӑ�X-�\��韓�TM)<*�坓!I[4e���Z���^m��W_`�)��z�%��I�gss�k=��Oz�� ��P83AJ9Hɧz���J���z}���Y��E@d�EV�'�Ս$�	��.�0qX"�T$�0�ŦT���xP_��Tb�_���D�Ҩ<yV�M�p>�?�GS��o�F������aV��cIc��|��[�J�>��������05/�V��y���7��&u@ �����G��!��a����p�Y��P� 	zy���tL�����#P��~-�0�k/K)V1w?P�_��Z��r�V+R���ǈ��<�DaEp{�Nw>�y�v�v��ym;2����e]o�4K�������i�Y�ax}�j,/�i�q��o�%�$a1��E��0���O*_"I}�|+	�9���e��ƍ���(KCM*�R���ϥ�G�{���D��8�-�+���"�	��
ڽ�y��Gi<����̗T~&�"�H�ԉ�^��B�MTaOp��L�����u���RǓ�Fp�2i5�9��{���`��4H����;.����)/!zh<�O��v�/W�$]� Pŧ�!��y���I��t���L�#��tXt%�v��A�Ճ��B�U�z��XU_�>F�eN�ya�S��
2���"SsY��5�3��~$g�ۀ��`(ͅ0�p.^�ܪ�ǼV�x��@�v��A�F+��mT3ݜ�3��8.r�ٝ����R�J���ѡ�+@v�*�8�W�.-�8k��p�lPT�?:����F�9*�\�K�Y����/Y^�1{K���<�`p /U�k�\n}nEAĊHn�[�|`�"����>��^ʽ�:8C�������@<�˜�!��ɮRjI�U�����t�N�BISbk5�Yf<��gڄx�"�`�EWS1Ҁ�P��5 �_���n��8OX�G ����(� _9	�'G�+ʄ�
d'c*h`�W�p��o(42w�Z<�c�U�G	��i����p#�۪m4O�)���`���@_ӕ�^�	�܏�A���ڜ�����\~��R�_����n�W*�C�l��I�ΖU�9ߗ��z�lP���#|,Lב��4D�;t�B"IbH�[�kek|!:'E԰���Q���[�+�Ko�x0ch��'�0F��`�t�6�P���
\�ѳkqI
,��������
�{��!R��A��:ʳ7�*����1}ˎ_�#�����~Y�~W<�+"v�� I,4�� M�zd��2H9C�t�T6���:ߊ�Mw�]���	��[�̑�UD��M��5?ou|Lq���+�^��,��?����oO�_7�/�u���W��һgoڤi�.DK��Fx$a\��M�9x�"!�[�.�H��&elV��w��[� ot��#2��f��[���[�I��xZ�"����{�FB�)$ �M���������g��+�4L9xt�48�J�����0�ur�Jv�KYTl���Խ9�Nu����$����Y��mp�m("C֮b>��P��+�D�|Sy�AݖP�z��g���=����j��
va4�z��q<�����ۗ�۳O%��T� ;,�z�e��s����77p���;�tx;�N�p���h���⊡��b����jE�t�Oy�������� j���$n����V+L�(�.L<R�-���@���)͢�@�)n(Cw�*�]����PmT,˿D')|Pk��f�:~ə�
�����4�1�8S��榧w�e@���=ܠ��̈�'l�� �ͱ�H��vJ�Z����e8���Dv��J]�����6b5�����#(��X��N����L�|���-z�~p|�R2�e���U
6u��9��Tkaa����bi��tb�"e���1v)�&�S������l�?l���o���41#���Zo�3s��	)�%hx��H,�� �����(L:6{��r"[1����������<ҋ�#��ɕΟ�Ct�C�PT��1��`|�͈
-�?6��-x*)����B���x>a'�L��v�q�v��Ig���ѳ��ɰ��p�����ߏ�{C�\���h5zI�!���������~��%��So�@}�au��zU����tˮ������ A,80�>�&K��Z����S�uc���a�z��A��{�a�w����:e�G8Q튐�
Y>6���q纷J?i#�/�9��gv[))��c���Ze/AҸM�!��.�4�5��ĺ񸎦�y��K�lr�R�t�b�q����1ؤew�zaza��܇���?����&gEA`ew�-�(t�\�$ZH,+[W�b�rP�6���� �-`T C���m��<(&^�l�񍗃Gq�C��>@�c�A!��xg#RQ��ꗺ���j��l%�Aۊ�[\<�$۠H��^�jH�s�2:Q�4�d�׆�����II:<�W��7��9�d�
��0 �*�	N�q,�	P��o"iY����I*��Q��ޣ���UG��Q����_��<h�cei��ĉ�݌�~K!�7���	)�;A�� �Г�'6rz��游1�BƇ.s�b�H�v^��U���5���A!"����^��-Ϯ4/�ghT2���oq�u\vX�h�����OSp!-�P6c:�
/ �����'�%R:�=�[LF0�s�ٯ�Gt�����{��,5&Ȑ N;ATO�˄6�7���^zL7���f~�[m\��"4���F����3��Jq�� ����g���$Ag3��~t�Rǌ�!�IE��~r����y���>�[ahC٨y��O��P�V�$qϓ��ɟj ><^��j��t#'��5ӈ;�s��式ߛt�����#�������X;@a^�]�Fg������mPԷ�;q�Gt��W�@S�֚�X�j���'�t?��ыڈѣ`��ei�82��� �����H\��/�r����97e֚ڳZ������I���m�0*���%���C-����C�{�X��e��(�6���ϔ��|�N\vjA�����zv����~��f�G8��/y��O�M���t]�a���ߘ;�2%��G�o�5��V�U_�T�m(�zSخ߳��&�BP%"ި2੼��e���s���X�é����Xˑߤ7���d절�<bl_�<"��ǯ `B�����3�����>��ݷ�*D��z�%��C[5r'fM��G1I݈To�Txȭ��>�6�e��1�(�t�i��v�I���a%��j��̓;�����< �{�Ͼ$�a�Y7�&�����i)�F�8�"�sa��BiG���d�LU�!D��\h��E�8O�����H�k���^�E���3��5��R�]
���w-�T���7��3�m�┾օ�}J���qY����~<ג��{�{?&��g�ݴ��^׬�GGEH����4�|�4��rG)��4f^�6=�MdJ����)������6�]�nHF���yN�[��m���)r�|��1�b~�aD[�ɔS�a�� �iC�|�ɪ�ef�Bu��M���j}��K���]�z��mȋ���l_o��VZo{I��v�6��!hN5���}�k8�ت��v��#gA��jD�o?����+CE�����u�in)x�x�U�5��4�C����
7�~�RB�A�)i� jtj�|�T��_�Oj9�4����aؤNS�0ڄ�W+B���|������Z�xܕ�R5%�n����fS�CY�?���e)L�ȋ!6�#�%���f����i��Xr� =
��?�B����u��kf��ILh�~��!������q~aة!9�&�� +!�P��юK�yIu�qFm�ο��Q����x�#$�D/4��<�r��E�Թϝ������3���K�F����B�B��ix	��K�	�k)���T#QY�ܱ��b.�2�a �F�)#*� r��F^��m��c�zbe��x��OakN�^s܎�C�<d������m �ڍ���U�V!y���U�?�Y*d"��h�di�PaI�ؓICO�f�k$�����Ɯ���d{����\�j1�$�M��'|�I~F;
�(&p�i#A�M7=��%cF2�V cD��Z8��u�=��[x���v��?nMM���� �p[3E$d��UA��TF�_T�cS,��.���@�R�r���t���?�������vg�K%1Sj���\����m֠� P�x ��gT�H�7�����g�I	�p�;[�׍�L�������T63����«����7�O2C��"�jރ�L�+`����V�HȾ��b��x}�g!E>��v�����{��:�}��ݘ�Da��U�������T��#S���X¯0��.Gwt�Wr��/���X�v����8��=�0أ䴖2����*�#qܻ�R}��xF�RK�7G��l8��U��=ʄbn������<q�!~���ǡ>�8������G�S�;����F75������D���g����,���z��sQ�g��V���c������� ��"?:����Y:<���0�@��N���(��0)�.UZ�����]�D*��Č��\�E�R��lG�n;�N_"�o��J� |f�蘛lm94��e#��5�O���e�Ĵ��i-b �/e�%�G�o��t�{�.5�\*���w��)���UҾ{5�+i;��v �s#�^��e��*�|�+e��"��I�SL�U�������׃�<qv���	�X{�K:[�*Յ�%��K]RcI��x��3�<QÓV�7,�1K��دS�W�2e^�D"���,+@I�Ӱ��3���I���@�]�e��w�[�NpΧ����;�V��C�ڛ�����J����]Ν�a��A,
�k��6�����j��$�/>Y4}���'j��D)�H��H���2��!����¢o�N� �)��u�� w����ȋ�?�ʄ�wq��Mɷ��DC����NTtXٍ��������[�+�Mm����	1bb�p�/���OE�B�F
#9 b'-�}j*w\J��mE�@z��:�D�}F����C����-��"\ݙ�6Θ����N�/P���(W�)�9W���i	����z=;y}��*�ő��ʻÑ<�4�4Zjܴ>"�*-jLE�0�kf~L)��~v�\�uF����w5�
A��:��S�#�����(f����<������#�6��Y z`�:/I7 }�^��ਁn��Y��Wu����7��D�k@�Ll߹�l���}'�J�v���b0��]��oAEe���X/y:�,��Hc*�y�l���;�U����8�;�x��B"B�.8�#ٗ��*��H��A��*îۮ�Gm�i!����Z�݂�l}p�>a��;����ܫ7o��BQa�{!���j�_��:KT�L��G�ٯ�%�ї�3ɚ�� ��h����tx4=щ*m=T�t3��Z��/�P�za�4f���}9�R1\Y��H�����d���4����ֈ8�\� mB}0Ǡv�u����xz��x��ަ��e�:*��x��/`��hT��H��f�5�n@"#�JG�U��Phr+:�X��PV���彵��z28=lt����/)�J3Rm�
k,Qj�W1utM���R��yեK@�7�tɑT�T P�N�"S?�^C���ܲ:4�??߆9�>���ϱ�0��m{J�9T%��%ԡCc��t���!���X����MH��RY�bKy�#?T�E��.��Ҁjps�G,��"%��b���
 %YL���_d$W���#1���g�A3|IcM�:v��]�LwC�I<��Ô1X4�~���>ρ�e���H�5�j	i9�����'��J;�J��e�B秖��D4.x�O�}4���X�����ؐ�X?�z�#Pƥ�M�%����hUzm�Dg���%ߚbѴ�x�?���w£��<#���3�i�O���Ȭً"�B�Eq�*D��bz�1��j�ހ�@�<<�f����M��T��QA�pHv��
{P&��AC-t����f�(,�o<�0�ʊ�5��~;��kS,�C�j���
�r��Kj�r�:lZ�V�m��`�;�,
�@H���{�A��r�G|Sx��1xU�>2�/Hl�+�y.�_�Dd��X��Ku����P��G���I�B"3����f�WͲQ[�qԑ�lV&�3�N��ɑW9���k�hYn�~��ö-F��$-m<�<�A���\�V�b߆����p����7!�4O����:�#>a����[��0�,��4Zg��YI7�9"���v#���o2^����h=�8?�qj�j��
���p���ʼ�ޅ��Q���Ղcacxd���	�b�=�yP�(�L1X��:c��������j������XA��X�.��_��1�T�|5#8¡*У~9�u�`�3<� ����ܥl	g��*�E�:_kn�_8u$d� x6����0|6��f������ɯ��i�-�%�^�� ��EPe~{=�s�������"h�7�I��$Z�6�I�����������V�W����"v� ]d�E�2��.��HH�7��g.����vK��9���I��j�#v�4�+9�H_���^C�
�������	�CRr�5���c7�=����C%]奂i��R�ʳ���ּ>#�����p��_O�_����D�Wq��C�cIE��x;*;�~`!�փ�9�0�K^=���''����jڜ�D;��0K��LƤ��NdkZ�7���T#c~&LE�߳s��^b��r��]��=�k������s��~o&� St��o�[NKq ������x��k)1�k�o3@�i!;!)�-j&M/+�΄fb�M����DtE
�R,Ʋ�֒�WG����F��&��:��	m�ia�9]D?�p��U��8�{\B4|UVV��Zv̈́���kFQ�����C�`W��;9V;s�H�CVy__*g �5h\�0� �L��i��T�f��U�|wn��z��5��ч�;rX���$�,�o���k��������7�����?b{��-bq6���h�����y2�3����rn����������N�D�V&-=�-F
��p��h���r�ds25U�GxW�_ցo5��[1U�:@�a��O(�7�F&�X).`=��&�pO��!_���yb�.l/9��|��CKx}]^x'��VF��/�2�8��i�c yEo��)ʅ�A�� hK�Z���>a�.6�p���F���iB<'��M�suo:h�as��M���6�)������5;���Oa�$1af�F��!UI�A8�A��<��<���6[��^y�!�xBܻ��F��BӦ���,�����Δ��j�����;#paԚd���<�x��|��#��$y-S��e������7�s������i���z�N]����26���/ �A��� E�;��3�=��.>^����˼�t�" �$ 9�R"��Y�ƩGY�4	�	wGn�y?��#�l��lx�x��W�r]Χ_Ԣ���Ԫ0�+)y}��V�Ƶ�$8�/ȷ'�VXyz��s�0@�p����7��;�V`�H���PJd1�ͥ�@CQ�STHC�v����݆���I���B!��=�5[F������`3�#���2؎�jn`��{�w�����i���b���큲O�R��Ъ%�"�n�<�Ovz+���.�d���Q�M%I���ޓ?[M 8z�ἣˏ�ŀJ�q��BK?ѻNuFzߞ��qQaQw��a��>�Gm�{���g������}��ܞǻ��$=S��z�,mW�Ҁ�AWDz�~��҉��!`���7�����?�(|7��ʶ����6��VC�`�N�?��	��Ei���L+(����d��M�|ħ�����O�;6�T}���Pe5�f�E��c�W'�������N��pX�Lo�/K�����&C�s��GO�76�0�������ߠH��N!i!�u�q�0���=�.W�m��@ք��vP���n9�7b\���i�s?��J�bk��W����p��$B�m"ҁ{�rH�k~�P��2l;�����$�e\���fo��4��]񘘟�ȟG>P����l�$Ȋ��Jsb��IR���8�3+G2sa�,ua�*�07�(����4���w#�;���'��E���^��?𺖈M��k0W�y?�{��S�
58����#|�Y�2kU��WC\wM��	
2�fh�c6A���*VJ�
��
���,�)(i+�7�[�Bx��%��, f�$��h큨��T�ݿyZ9ݸ�P���n sr�|�墳�WD�x+8�76��qs����m˛�p������`\�+�1���� R�#��P�yyqܚY��]���1qO9	ޅ������a��)
<�Y`���VY9�up.���ٖ�G�I����aT.@����@I��4d܀)t�J<�]��S k�;�	@&���R%�	�֋�+�R��]i�D�H�Ha�Y0mk���/m���^�?aQ2cfv~%%i{��F'$�)|���pUVj%B-�q�?��YOD��I</�����*�cK9}o��t���3��~k�bw��V�1w��TǮ@�@���ȼ �lWɊ!�\��/��l�a�}T�ÿ���*�Vⓣ����i�%���V�FԌ���o6���.��;��z\�b���k+m
� ���$gǳF����xt/M8�Q�ۺe1R��V0�X=��-��,aC��#�9��X�k�|��agb��0y�X�<@Ҍ���(�������Ԛl&p�ށ���z�Η:i�3V>��RkV��U�[� ��s#���γ��$���?�T
�G��C#?hĢL�~��*.�;"-�`Ԟtێ���\+���hw`E�<���E�?���?qF�Ǟ�BL�"�o�A��j�6XL��'	9<K	��}�mS8hYg���e�N��&Kc���������E�x��M?T��MN��f#C�x-�,b�a�l��,�8��H�uS�g*@-1$�qa�r`&/L���em@Τ�!!��mǫ��X"wU��xq;ګ�"7Q���R|u�VsT�mb��%3d�	�R��yF�q�l��Y."�M�V!�|�X=W�0x�s���琻��¶�G�/5e��l�t�2�Y�b+�5u�k\�
2���+��S��P�ZM����ce@�G|�q8Ke؂i�������S��M@�g��1��֊�ܓ�^8��!I�O�7J87�ü�� q�E&5�5
��,��8L�3�����G�}R��Y��4H~f��v7��p2������&���W/���ii���S��4*
{�� "ol�b6*�� ׭L*��;���HT�F��K4Kʝ��N8nD�WI��� :E��S3tt�����4Ɛ�II2�^�wFߪ��F��Oʻ��1>������M����x��p���ai�c��K�S,� \6^ݑ�_�3{�]>q�����K����M[}�i�����č���@6�������s�},
2o��!'}�;OD=6�Q+G��k�㣸���79��������&����K�cC���a�d/����#��q�4��r;i�6&�P���)G&���o�����݅�������%T;�\�����P�Uh4x��R؋0i��Z{8�\S$G��f���(!�1�P�N7�
���-rh�SP�4�P�ʌv�����WVgx�[�<��N�ryq��P4��h=��Iv6��pq9�e�'������O8�N�o�����2eH�m�(s�2 ������>�k$�Z���׆����~#t�j���r��gʳ�=|ʯJeB�©�#$'{l@}c�4�Q��.X�P�,�#�f�O�|kع�J�kņ�b�#�,�VY����D)Rw9	f�a�����Ǌ\'>���w'���$��͡ ��Dv4{�9f5���n�y3�4��r��M�W�٥.[I;��?�V�֞^�F��"�_�\�>#@������R�k;f�3���?~t3��Pn�6�$f��F f�E�m���	[�#HJħ1ȡ��� lHw�@zݭ�̍�2�����ԧ���Ã8n�^���&��O�1�PU=^�)3^�%�FM�ܨĸ|sI��f䁵����m@vJ|�X�|��&Z�+������qf&��)��`��K�ӈ������6��h:G�#޺���#��������\�Ѐ�,vE�����N�<֋���5�S@����oN�i7X0���c���ToNʛ=��=�_�r�㻉nTQ��D��H#0�:�^x��J-����b(�����������M;����}ս
�6P��8:�͐rgfAa�=ͷu�?����!�s�[������'�a��L�Xغ�&"nJ�Ȓ�"���_L���o���mz�X��k�E��l�� :q���5џif"�C��VFs��Ҏk���sx��8�f���U�rD�^~*V+}��,����ɑ�� e�>3�+rZ�7k|\�����"��5hB���k�羮g�5 �Ze��7��o ڣ��+#\]�:� �~E:��S!�nbOlf���@�0(k�c�[ɍ��?y�;c��v��S�(���x�<��0������[]��������(�ݕ8�O�CU@�뤱�GF��U�֌&�k���!h���U�HkS�?_�Oy��Z�	�M�0�93���=�b�����(pt�d�Ns��X���3����Uo����x$���,���;�vO2�ǭw�{u? �W%���ޮ���q�/&"!��F+����i<��^N�������yu�e��3n��bicDeh7{2ۑ
ӱF�="�r�!��lYxTj�e�l�27.�KVX&��/���1��	ײ��'a0o�U�P�{8�V�2�M"_���ɗ�\ݦo�|�O���8n�q a�}��[ ��?�0��Z ���ù���Ҋӟ�v�P:��Ԡ�s�̑'�6��&�����";�3�LX`�]�	�5� ���UN;`�\�u�"y"�����MVd�]
iw���y��-�$.)&�)��@�S��z�/<��t3���O�I�� nL��o�`���D���]~x!����~'�d�P�w��0�g|@�J(��gn`^7��I֣�w��%�G�g�����n���0��(�y�SӁyrT�3H���܁`��9���x�`j�C�i5S![P#>kK�oX�G�����b(��^nB��m���h���)o����Ta�h�ě���5�PqT�6��D���ِh%�M���F��`�X(����>>��i����8�`�T3�����<�^4D�SQ�-��S�G��Y�&mB�;�ˤ�������n_R5�:��
�	'ٽ:"�`�Z��M�}s�㳩�E:����]��AdZQ(L	��ݖԩ��f�ſSd�r��ڛڷ�$�H�q_���V���H w�7����v�+������/�(�r]�Fڀ2����ո�Xjf�h