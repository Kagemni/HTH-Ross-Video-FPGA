��/  �F�o�~��csT@�e�u@�� ���c�;s��H���W�}m�5|�p���˖�p0�q�����-g��zI��N:ϛ�+x/�Ps;I�r8'���!\��E���5��32� ;��U5�Оa*ʺ�b�9M����V�ʥD��/�q�2큑��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�UtK��^�)A���Q���=�.m[�F|��]C�9o���m����T��i���`3��.uFh!%�S)|cph$��ڞكRy�4��Ӌ%ǖ� ��	pv�.����D>g.��?��8�������!ʌ�r#�ȇ��
�<D�v�$ͯ�=�Ŧ/��l�Ϻs���ؾ��@��;�Ǣ������������ج�@L~���/��dU�����S%K�xW/�E��ĉX{.�X=�? ����;3�J�-%��"9-�x%i�tb�ʽ	|����:��U��D����<���;M����h<c��P0�܃���
G�v��B�7G�j������L�����D��Y���e��!rF��G�x?���f$��s��S��	��^�J6RD��Gd��t»�����Cx��dib���9W@��e�c
ӊ����!Y�w(�	�*<��7?^��S���$�d<1�t&�;J)�j�|iv�ΘV�I0UU=6o4���lU��^O_ŖhK�<��C�q�z�L�m���>?<��F�lW::�r�5Ob���,Kt�L��A��x��}�݂Ҋ�뉝�'`@J�h���<��ĺk ���* ��u��������UI�'e��%�jsO䤯�D���7}����+�a$4�T�׏E�����6J��z_b�j#�^��GN!�l�2պ4�~�"<;��V�DGBh��LF'E���o��Z��+�ж"�oC;(x��A��}z��
7q�d�O�6BAf^C[����Y�~���ֻ���:��2�u�IP�# ��tT��hR��*E^ea�b�	�F�S°
����x�[Oq��`��Oc����ڻ\%���ֆr�WD5 Q�y�#�3��^m��T�C��8A�՝��׶W�]�B9P�H�"ƙx���ŏ����0)�{'KtD��ˉT���|-�Ũ�EM\�m��/�4�ڑ2WK��+�@�����m�5Ԥd�{K6�lr���;�q���j��1�����20͎Fw ;Q�=�(��Ȏ�.��YX�@��ݳ�<�l%��ۋN������@,.P�G�Gw��P=+�-��%D���CV�qCIG�����i8�k`=�C�x�:��G�פ� +����־p���QQ���E�I~�ې�F�l%t�E7��]�}j�.���icW����$�p�Z9Dd��R �6#aL��	�*��O[��6.���RY�~�	4�{vk�` r86�ʑ��V�ϫ�r�<tl̹�.�6��A�:��5}UǨ�D ���HK�ZY����x�}�g�T2�M��.{+c��gi�wq�j��+��;�a�@�*�S$�e����9O��_ f�����z<���'��5C�I]�ip��~����;=��l�z�jߜU^4�19f��<7#�p������a�C߮f&>�k 8��"�W<��R�Fv���܍�G�L��>GE���Piή:���E"�B�_^����?�z��|��>�>|�f5_�+�U��t>�\˼DT�2��I]8=�[�ԏ
� �Dfǽ.|+D�E.A�����Z?�>����.ئ3=�˵O� ��7�A���J�Y3����i]��N���	���W˪�#I!H�^o�P�B�")x�&~~#ӅB�D0E[	�r�7��P�B�"�C�z>4m�rBm=s�:�_&u��]8B�O�%���hV�O���_��tw�ia�����#�l�T
�A4Y$�r9s�Y|/�c�L�2F�h�����T^����kp#3�H0h�^I���o�����{���p�ǥ��F��0eA9�Ua�}���D����ʊ� ���N����.�.%�uk�8��6���WK>N��@�q�]�)����}�K��&ݎp�	멿k����]��ʿ�t��2=c�ݷ�Y�� ������NX�1�̘lXe��P�Ֆ��ҷ�:e9����?��Gd2��!AE��L�u���h���%�a������=���K&�o��k'���:�3� �,�]M�*)�49���D$u�R�B x<f��*�919t;�I����b��O�k1�׹,@W-�7�6�招�E|�g#q�qXk�y��m3Lq��,wM#YV4���a⫹��rد������5�8�lS,l����m�w3ک�&�cRSG`��*�pl`¸��.���9 ���"�I�����$"�78����h�q�	e�a��G큊+T��V��HVWA{9aќ���7��y�uJm�5��ښ=��PY�(�,�	y1{:u?�Y��׫�K��#�Ik�#��,s4L	�əB���u�{��\�Z��BQ"β��^���`L��Ӻ��3�]f �m��+2ɇ�\�˼	ʹ�!>�����W|*S/x�_��i��w: ��i�1�7��q�zJ�0��،ɼY"�֒���r�����J�~V��퍓��$gJ��q:�־"�*C���f�6����rP=��Q4z+�X�@
��m6ԅ�e~ݕI@�G�\O�PBd��|��G�4�th:'0@��y�Y�L�&GC4&� �.`%��U�P�ha��
��&Ms���gU%���II+'u��,ǫ�R��̉�.�ժ���F��&���o ���=y0�n�BD�/)�#�U��na���;�DV~�m=��S�����I;��l�ߓ��#�g�n��);�P!�G�Ȯ��נ��]���x�B?V��7��$4ʩ����L`����b09�� 7rgB�R�Sz���4D�����P.���0�=js�����*���{3�5d{P��u`�?xe�`.Ҳ~NO���
R��������1�v ��>c�y(
hvW��X�zA��D~!���;�z�� �3șY��N�鉌�_�����K�X�$Ή]�;Fo�͙^���l���7���_ih[wF��AQ\��;9�qt-;3?x�[����5�(;���	XS�P}P�S���r׾,��8=ծ�E����Q,b���c4�u��.+k&�YFk;��ꞟ�y�����9^�X'���%S 6���I�9���3�"-5 �'�h9��а$(������h��g�k���`��v�����
^��$�vɖ�����
��`H3[��J��d�](���|-|*wnnF�:�)��[���k�+Ϳ��I�C�L�"�)&f�ѹ>\���)���q=�.�.������B�̨�Xj�i����`�#?%��e�vV�$sp��!+^M��� !xӯ�	?�L4���q�N�Z�A�',����Y���+��".͙�}�z^�,m.���z:���&��qM������o�֬vQ�J�>�7F�G+��C����m�������X2�g9��/˺�V��F�Z}	���H�.y�&�F&�-��R�8��>�;��s���p��M�nCǯ��jW�k�o�$2e��n�n��}>���UC4�-���ZdHƙ.��$ˮ�����t��WM����d��uV��4�����ߘs�����y41�L�!���s�ǘ/$v�ȡ�%�S6ot�nG��@��:�q<6$�e�����8n���'�\z�4�;%gB�\{����.��Y�H
�H��|�ff�q'D1?�<��H�1����a4+HبQ}=���(�� ����rsBvS�P�쏆Ox�~�턭-��r��Sú,g�@����ȭ� R�izr���S��Ꝉ؊�+��.%�\�{^�e_4�9�mo���^�!�v���cıO���~d�G-<����WkOC�3b{�u���AM���`^�u�lLi'���_�3ah�6P���!fp��Y��Pu�F(m�C0��������7h�L���e�#�t�3#w0K3V�N��?�~K�������� �jӗ���?���R)O�e��G߳����'?'g7�wW�LCf�Q�`"��5!%5��d�� �2t��~�r��ҔƵ�\�JY	�)u�P�&cv��ӣ���Mb�X�ͣOD��_q��J 5��3��V�ZQ�a�RE���-pGJ]''��́1���,i�����'���@P8j=�F�mi;f�Q��ÅT�xe��$�x��V}`���_53����<�ě�S��_ҋ���<�Yg�[�w����,J�ͷm���qp���ju��`W���a�U}��!��{(��vQl4�K2�U�vd"I��'���m6��d�H�;���H\ ��)l�*�����dn~@��*��`ݣ�u@P���{V�!	(��?_ؗ)hS��*䅦���s<T2�,S]����D񛤐$7a�����İ�	Ԕ)�K�p�{���)����nW���8x5�s�o"I5kа��w���5��G,gM�XA���\������+���
�B���r��_;3;�x�rcz��9��̗���M�ퟒ���;�w��t^��%XX�A�G��]+��1@@����~F����YP�\����8���p��`�p/�L���3b���P�o9�:���e�֫/l���4�Y�6 �_�H�,ތOk�����Bl��"v��b?�<�����y�m�8�m|��R^wݥY��`��1�)5�!�2Ml:��Є��8�$"18����'��1�5����Я��/���EC4jVT��^���z�3�4�6��=�|�w�����X:\.�y�u� �3�e$�չZ?2�:�@IBB��k�
D�|�j��OI�X�K��<���M�w�0g�Z	�#��WB���l���|�mf���2��(�*mZ��J�k�1��Њ�)7�,�z8!��}^�Je2���O�3Dx!#E���U� ���G�`�5��L\�s����)k���y�PA��ׇy	�>��O`��RJw�g����X���^	(DLx������uqjPrZ�O$���K��p�~|���ˏ\!�6S���!��=�ӓ���������`���������yo����e��oT|�
\Tzb��\	[�>�!B_\9��QI�E�}t�
�8}�3ൠ(H���:bX(G�J�5?���"�FY�`ѱn���1~g){���onpXMA���$7D�����ԣ>��j��()�e������{u� �p�x��&M��hbY��2�����f�-�z��l�1&�c�%������<+h��T�(��g�+˪_a�S��#�8�`K��*w��o��ą�|R?y;�/h�O�?*f'�5@�8_x؋��Y��h�gm���լw���S�^�L��!��Q���KZK�`��3n��n�ꍄԎ���/����әE���y���0�J���&�l����yت,�
�}bs�&���-�B�S��O��_�s=�B���t���k��J��#z�R`�<�QW���?g��[%h^�}6�q'Bª���v����kK�Z�!�	˲DG���?>��n�[��a/��s+Ǡ�tt������->�{d�*ZJ��Ӆ�-�ZA��`Y�'�ª3��F��蛜 ���n��M#�ǌg�30��6� ��g���K�{	��OwYl) I+��ʀwm���Up������>�A=nQ.��q#]ŉ�'���}W��tn�i{'�:���b�����'����2��FM��-j	�X�ӽãOy?|��"��j
�����X��F㝾P��������b�����I��Xl|Y�P�y<�u߸�w�h�g_s@���:���uaijލ|B~"6����8�����;!;̨�k���)g�^�@�e��pz>��x��_�`Z�rZ���o�Q�Gl�9o�q��2�$�󑇞%s��4�.3�)��
C�=VE��A[4�-QH�e3 �>����]?g#���#���cyr!�����XV�U�k��7����îQz�
B�#:a$��Ҁ�� O\�,�a"w����8�)>��oR�L�m݃A��^�:hw�um%&bK��MιQ>s?A��P3�}����G��M�B�Ǽ6�*xj��K��>iXt�X,���O]���G�9�yN�M�lo.�]M�Y����yu6n0�e����Zsl��ⴢ���eQ6�te�@��7yN� �S�|w�����3��0sғ6�R�q\�îx�ʈ�DP��yT���/�go��ʉ�0 ���,7z��,���cըM�]^�`8z)q��gk-�~��hr=�����\��r0	m i �V���@.��DEyRZx�M���§��r�Ǭ]����0���o�3����b�yPի|g.�9�g��4�?T�S�7~
o�F�"�̤�mA�<B�w�d�I佱h"�$����(�e���~��8��J�4H*Ea��F��b�{r�=/�(������Q
|Y�˭B�+@�\E/���z̖�h����Xb>���^J���'aO��N9 ����m_&�����j��R��n�uǒ�ݕ��/D17.��f�~���nԶG\�P�h
E	�d��#��$��uO=_��E6t#$s8��
��
�◳n���˿�=X�D�r�!W��B��=��L���hA�e���م`s�?��Zsu�P��ެ��%�0�"�;��ҹ�9�ᤃ�zN�t���kE�j�Y�qCb iO�ˣO��g%��O1��0䬝Vq�I��*�<����oĆ��E�|�W]�q�6�4��M*��m4흦;��7�V��~���/t�t!@6�c�{���֯�I��}���j�
"a!�B��6���y
)���ښ�I�����|��Z���f�Zć�����O� �}x�0�� ���ؤ��R�\IQ@��Q�\�_�8-�E4�~�Xx=����!�	0G��-�ڧB�tGDdPǅ�+�6W��\����t�����k!��²�d,����H�o��8!V���z�us��rU��7�V7����;B/��c ����$��#T��g��)GѪ��*EbB��@���͒��P� �vf�i1���ĺ��"�|?���vC2_ɵ�ƣ�k�APlγ�:mӸ�8F��1'��,����ؐ `8�yg��`��"�9�_�>� ��/�����q��G�cjD���6N�*͋k)<ܵ&��r"%-�e(*:���Y����v�HQ�p���㤥l�M�1�|�ᤸ5���΍a����b���/X�U5M	ev�P���2L}���5������C�--�j3�t�o��1�f�}`Q�/��:�{�C,5aA��>��_��^Eg\�Fϛ%XK��<��>��y�{Oc1l��B}���*,��e1!��'�3/��_
�Wd`�V>/�H%/�/�/�X����W�ހ�ހ�}~�Ǽ�n-�kh��B� �`g[��3�u_���2j\X*��j.)}�#�]U}�R�/�W���뚃۽�˗s5vk��!!��-{u\� ��r���ƶH�/���zWH���W4x������Y``"nPq��U/��8C��ٮ�';�A9W/I�}���?;�x��n��Z��y݄+�I�1m�۳�S%@o�S��.]�]P>%p����p�J����u�N�ί%
��<F�W���8*>�1�F@�o�K�����,�_y;�>Fi+Pϗ�?�l�X<��] �3Έ+�k�{~-/���q�� ӵ	^����>/OIXb6h����S{�H��ce�x1^5~�&�7�]�:�L�ٵm̦G�s+�l�n����s���}�ږ�����S�7�f���D�M��
��\�x�Es�$x�Z3��^\�$�b*�E���$5��������7���e�x��jp��dY 4��}5��<�Y��RB�k�L��f;�}SoV��&13��'� �^|,'y�V���hO/Ȏ�Hp���^���'KWA(��W�w�@�ۯU��D5�ZE¶w�Z�f- Ky�`t(���oQ���L
�%����r�Rq�Dv�A⨘nD�ZS��O����@4�Ip�h�+�E�\X��5H@d8��<~�Z�l�2����{�uHSPz'����Kt��qL���1��~}m)hDPg��(��@+�蚷4��N'z�[�����\�h��"�)��.w`�O%��9����.�*G�$}5�H(e���N[�ƾ�5�Xľ�2xԙJ��2���W���z���aĩ ,�[����k���s��,C�#4�	ú��/(��8����{B';S��7<��O{G��1���6t�C�b]-�s�}|���'�F|�E�~}�I���!��/8Lr���Jۉ����5��W���]��uB��{Wtپ��.�ɓr�O�F���T۱r���>��sM�1��K�Si�A�\F�Gq�V�Hm�hܲ��B
�6���S['�>�����J���2VOy��Ƕ'�L,"������ϰ��u���%!Q��=TQ�MɊ���`0�����{*/u�#x��xm����%�1#c�I���8O���)>vn�X�>|(�];���	���Zʈ��S����U�j������Tt�r�Y�-�3��qZD`.n��jϒ1$�R�iNqwÚ�����?�����ڇOJ�| ���I9�����Ѩ*���
J��wD~�ۙW�O0iMݛ�/��_� <8�����?�MC�3�R%��ô��9�vr�5v�	q|�c�/�l�ot
lF����ĥ��-��q�Xj�Q%� i�p�Z)��!]݅����4����VS.���E���<"���}+��},�2��[
�&H7G|��~/��\��"���+<�T+8�������`��Ǉ��Ʋͼ��_�ގ���T�������uy0�uZkE��N�w~q��3��5�`K����>K˭��)�|�+ML�8��rgΧ�����%��_�U��k����������1�W���SE�F�����L�Gڑc�y�y\�F�k��7J���o��$>�e�eD�cA0YY�a��k�;-?Q��@�NN?�DR{�/TH'[s�R70&��J�E�θE���*T���TE;Y*�5G)"L�5v��l�R+�nA�彀�A]���>����.%��-�{��� �bm)��%-B�L]�	���d�?c���
;�er�ܧZV6Nެ�Zd���?9����@&P	p`�	Q�H�������^"p'nV��F�F�cè�(ね��o��.���l��DN�I�zlz��^�mu����AÎ
�gL��˭�U�%�q�7'9���$Ŗ2�{P���pq���⸖�!�������k�*�ÿz[s�2�Z�����)ه�0# ��]�r�/i�k�X�a�W6Ky7v�&7��ijTQ'Pm@��%*�y'�)���۴��uˡ�T+(�U;X�L�t(�&4�^�Kt�W/zp��L�m�}p5�(�L��
2��f:���p��D������'��L^�R̽l�~��;��ŝcCx���"���f��&,�9��~��S�;)�#b�Y��m��[�����+fxz<D��~����7���c�:�٭U��`h,A�*��Z��	�$�V�OW�,�Č7b*2W*V��P�!ѿ���g�_�~v���s���-l纨�Fz���?�"(�l�IHSTq�[eY����-�K�K�ӹ���w,vDJ�"V���K���A8NvX�)�(6=���
��@�/O?��K(�% BhV�x�$��i]-���TŤ��{sؾXǀDބ�B����P^yf(G�S/�9JfB��MG?�A�6=�9�젨�$�A�y)����Ādi���[�Kڙ����X�߹ �g��w/��No袯�!s���*��:���ޚ�X���$K���W���{_އ�b�8nK�+�i����YQ��#�]�.ō�it��K�� \�w��ϻ�%�����W8�Z����R�����)F��)��<��x�}z�쳩����4oq�~�5���Q���K�ғ� �}���6IfV�b�hi�;DpƏ�|�r��oQ��fF�;�F6�Ǒ���ՒĤ5�3�بu*� �M�����t���!/�8���b!�Ӎ�9]UV�v1̴��B�5��
��RP�2���S�^ǛV,��������[#�og�*%*X�� tڲ:d]2�P�I�
��#��y��U�",�jQ�F 1E���+�d�ס���AB>�j8�u�����\��}�PƢ��b��.s��k�Q:�;ϱ��*+޷��W'��Ǚ��ֲE��;�d�~v�^�M�di<���Ϯ+�N��6]��B�l�O\��^�}�fQ��Pcz��#P���K���'h9�~�9��˿���I���;Ӟ�!��(h������A~m-���u�p̫o�%�vn\;��u�ّyh�e�1r�	y[�]U��[l��i&œ�!��T�
�oyp�I 5k��-t���/b���~���v��Y���5+�0	�%�`���]"�LB�S�Ӂ�`	�8v���Q:�J�.�%�	�&OBxg<a��@v	��p�"��%�~��F�P$ŇE�:�8^�k�#��Z0�5��3|	W6��N6��L���U�qa��`m��aj'g�{qf~��>��u�c��h�ہ��2�B|I�X���5�H��<F1��챘:2(₉��\��Ӻ��v����l©���Q�3քL��^�|3p�!�J��aҜ.�!�]�/i.g1q��u$�l�VX���w��J���% �:���޶:��y�.�T��A�^Y�V�xk�H��[%W}T�99]@���ƛ�BZUd<?��"�P�U����TN�70!o�����Q�\2��P��:x&CR���rL�6�~"�	�0"�m48E��ql�v�����-�.��G�|ym(��i�~��3�y����z�}�����ı
Rd��~�����~]3N������x�w���</���45��Ӭ!n���n�m��L��	˯�{��_�0�l������c.�00�c!ŏ�ͣM1��)^�|�mW��	*3�C�l�u
 D�1=*Aƥj�6Qy3yrU��*��z먡v:�0��>a�Ψ�Q��M���P̖_7H� ��e]&cue|�u�+�!�wO��R�M�	��a���=4��q����EB�	��s��Z�z�Jt˟�鰽ْ�.�Lf�����5���9�x�խ�>N2��B]��;�MC�a��=�G����`�w%���*�R�iq�"p^���L�o:�APfR����&���I��Uψ�ˬ�)��Ap�!��`��q�4�����	?��Du�D�h�S��(�ш>|�c�rm�Z�c�"\�H�ݝ��oakM�y�q�������QB0:�h�����T(;A��'h/Ѧ����=?P~��I�,n"`|�X[�ѻHgyr��򍁝?�`A�
-@1���\O���=������ӘO��/���MWě|�}\�D�Lt 
�\�D��3z����\��B���Ԛ2��Z�8?O3Or9���_T����4���I)5{8!uFI��񕼑�<��Lc��o�1\�?MK(]����ΰ�DS,7j v{	끣��l��>u��۝dY�%]ޖQ
R];�����?
��R;�z�M�曅C�w �)|�7 �8�w8���7h"���&�W�����=�D&��Hj�1���k�(U1�4+����4@����w�0����ԓ %3��0/��s�_�NA����8�$c��(%�j�2z�� ì�iɤ�5T�Kv����ܹ������}�+-����*���^e��5l�	�$Yp	mv8�U�/����器��`�R�OV�ѬHW�8=30jVx�[���Zr�&x��W���%F7Nb2�/E�l`���aae�Nz��d�xy.,����([�����Db���4C�D͆IԿn��]?Q�F�)==�W��[�k�f>1~0��� �I�N�`6o!��+���4a����X��Y�/�]G��C*G�o(yЬ�Ƀ�X"~j@U4(�Ս�FjZ�} -Z�`��A���N�N����(�u����l?z<6A����u�]����|  �dM���|[�Njv�!�$�>6��}F���'�L�u�~�o�z���(��-��]|��qĜ���&�0�5���7/-�����q�L��)fC���u���֣O�Y�:������c�@�]o_� �# �oGB*�j�	<vW�U��=~��<���&+32q����q�������s��@���%�:�Z���Y����57=�
IdP�r�T|��8�����K B��l�7���"v�Q"�\-׼#��ׯr�gV��m@[�����.����0���t9��\�(d�5����<PR�u��v���A"�^�a��R5	&���p`e�JƬ��d#h���X�WX^���oW"�wY �EV���襷7N���\���˔qB&Gȇ�Ƶ,v		_f����_Q�$<B��%Ӄ���G�4�1~3|�����3�ܤ��T}��C � g�Z^<��n�y�O��u7�k������f_��$'��H���5�#�F�a����[�%h�����L���Z犅���]��˲��s"�|��(�Y�ߧ��"Q��ğ7N��%,���6�T��i���r�%������2eҗ ª��D��K�4���7D�X��n�T�;!��n1���-u$u��@5H�N6�X�!�>�<X�.Lwɺ�Q~+�wE�4~��#�lS��ǁ0T'�^�dv���}�G���Ro\0�|}��0�I�)�B�I�_r�oD�/�49C�ˆ��K
~�����o/����dC�H��[��1��'�d����pƆ�j���:����������� ��߿?"����`M�2*�0��V����jS��=zП��Ӄ#`N�{t�������3&	�V)"�^�.��PRګ��*������#^ [��W%�\���2��ܘ�x�=�:s�DtH�����{˰�"9�4�6?��S@ ���
5^�Lx�/�E&BDJP���`&��a�Y���aV}�@�}!`�+�~���Gi0Q��y�VlN��P�U���3X��"J�3��F�)��t�O..*mIq)UY��+�}]���^�J8���:�r��?tf��n$�5�x���n�Z1�|�J.Ԧ���>�o�@rG�CJ"[�Β��Q_����X@��� NeۄWkt�r�o!��*�����x%�1BE�؃o�3Yz8��p߈�c�i���쵀'F-1�qybVﬄ=q���G���j.�V>��}�|��yoY��O����z�d�*�i@�I�S�Rv� ^�U�?v)q��5�!��OQ
�W�?+,~�c�E�8�T�&9�,�!���q��觥�A�����~�&ٳ9%'��#/�t!�8�iQ,��Y/Yܨ��;��j�1�Ʒ�Ĩ�BWѮ"b3����CI��jjJb��(�NW?�뺘iR�I�Q�e��5�|b/2�e&×�X����mv�M�^!�L�4`�o7�I����%N5�8�	8-)e����$^�n�p�Y᜻8��յ��w���Y�~��>j�v�>�ʡ��Ņ���X�~�<�w1�J�:?x&j��ٯijO
��t�7��`��$�����ͫ�HnءC�g�k&#��\��b��#���B��}
�-}�T�͈5�'��2O��g�g�>¬�$ 6;�F3�j��fA��8�K�um�{��rlـ�)��ũ�t���9���C�)�A+�:�0�f��?e�z���C�r(ie)P>��^d�$�H��	̣`F%m�G|>?'ց�#�Q(R�65�T����f��~ONC��ݷ��@�2&�fvӣ$�G�gb1�A
�B���`�ؗ%F�QS��a?\��=�j�)](��s.-˱����N��O<��;�7��OUΣ�+����e��tɔ���.����?z��'p<�?��/�����<_?4�5�|�c�^�35���K��+���ߑ�������0��I�F=�1�4V��gX�R"o�c�N�v�w�yrύ�sd��dn2z���-�9���X�fY0�ߵ�"�](�$T�'}z�}�X�"GVȭL/"�Hy�u3�|�=����� �0�Ԧ�3���8x�	���f��}��0J��^�_�>ԋ�\W��dӳs���x��ؓ�]�a�:�q���EL"��$���j����>��G���Wm��L��GQ�m\�!;cD��?T��0g��d��|U2A�A��Po��ː��UOV���1��TxNN�刭���{���ʿ���gs�G�i�j��~LXX볘Ch��j��Iі�BR|5�uԒ,@�k`����Op_�i�TF��/a6t�ȫߜkrgz�>Me�.f�������Z�#�}\A�߭�E�ʶBqE�R/�FJ6 �M ���c@|�݇�>�cTL�ҕ�2`^w��Ɗ�F.y�����?����|\�$eu�B��.��~�:Q�5k-�u�w(]Z�\0 �[|S;�5QJ�6�,6f��z��Wi��#����G��E >�+X7Ĩ�j1��9d*�A�汢 //ՠU<y���à���ʶkӑ��d���|M|�B�3�c��Em��迹X�y�����E�S	W��$��f�W�0 lr[[�:��s�w}�@ΤS�2��U�(5:�
G���[.w��ۙ3mE��`F�">��X�Ap6P"ꂌ���*mC3�������*�w��[`�$�c�4�*�ꀖ���Yj����z=�*���!	eaCJ��V7O�K�U��x�oE��j�e��N���� ��^0�0�MU���)�@�+�����W�U4e;B!2��9��d+ciJ1]��&G@�=q;u� }v&M2�p*hz��oX�Y	1����r^�����v�x�O���]l�B�[�#�|��1��F��+��Q��&�i�q��%�ih�3�Ƭ�[@�vaZ���i(���a�q�rQ
�V:+1�̖���53�d[K�O2d�j<CڐM��j��n@sV�~
2G+�0o"�K�U%�B���<�c֊�ÞF=��pz��U3[��C/_�}w��˨��2o��x��~ ��ѦLb	�l)�9x�q�k���M�3�����Ϣ�UX�C���
#D�ġ�T�t�x4oGA�reZ'��O���4ܭZ�)��͏0:��FB��N��'�Np�Q\yi�G���f�s�_�����5[ӊZ1�N��ĚN�.�=�[@�3Q�~���9ъg�������Q��f���?˹hA���c<�*��h��I�C�������M�ח�qź���M��k��A{���̇;Q�8f���.��{SZ�b���H�\~qB)����DqDf��S3eD�l���_oaN� �a�=ٲ5k2/�>���
 UC��e��쌃h۪6�Ԩ��oaG|�c���W,��B����� ��CS��)'Q�T$Y��f�	>�(�=H�,�n�j�)�s�m:��Ӳ�={Kg�������v�g�rx;�����B���lƨq(�I\�!7d�Ht!����ؾl�3�p��>�����o����h����i��rAL8ؐ*���4��|;��MOZ��E�$��6���lilQV<�����X�࣯�|��aq"����T��D P��#O�'��\;�Z��V�)S�CO'�� FόA��
�uWt�R{gkS�#3U��ռ�_T��f[�lҎ%��?���gm�&��}"����s%��R�$<0�a���m5���!����ƥ���I�\P�V��zJ��SK��U7bTuk����.�3@y��V�?�-�j���/z�'�A�#3���FTL��~k�i�77PV�Z��$(b�z
ϳ�F�+���I<TL���lh*�h~�+�p��>�&_r�{Qk�E\�%�*_P69x���i���jޝ�ށ_���@��/�
��SY);��ǃF=��N+�<c����m�f2�:\P��:0�!c�;1���_�C���eDiS�s���O�,�r��ۂ������Q��`!�n��hnK���as����}�D74�Mi�B��==��S�
�@-V`��5Pץ����;�,;�<���ZH�ΞQ�9px��4��S?����BNG�f�-z���6��O�e�7^B��fa�=� 9K�����{U�B*�� ��e1�L�g���"q���D���nOD�킙e���/���D����V0Bh���~	��n���6�yjT���X������qvKU�I�rWy�#���
Ǡ��5mm�(���Zdd��R�#>��������lIm��H���1�l���C�I>��?&���b��,��&�X���e-�O��r������;:��U�|@p�R$(.HMe��о����Tk82[�h����j�՝#���}SrRJ��d˽a���L���i���;Y���7��ڝ�/�Оւ�R���Y�ȳq�^\�&x�j��"��)[oԧ¦��[�I�����7��b�O��ԉ�oWݰ*AxR�ٰ��,�|tњ��禮�}�ւ� ��/k������l��#4�s_S�Wz9������=9ڇ��C�BS����I�P�M#�7��u�/�s`�:O%
y9�ITP��
*��X!^�Sjt���^9C/\����#�����Df��Y[�+]%��m5r���O��O+Z0����ޒ�>V�E~���]����+	T�(u�㜕�C]t���=ѯ�V�]�'�։�~�r�����\ɾ,|��0�����G��Z�]'�lC�X�M돔k�Zk�(�����@>�k�^����;���8(U"�� �4��]�������~/���צ�F���z}e�����e��A�X��H� &�,JJ�_C;�G�<7�8����٣s|��D7Ҏ��1�b�n���v(½��W;���4�����TfQ�光��r]��E$��F���d9� �τ�̏���Z���V¯�9���x��j���L%)��[3����5��Z} ����B�<�>v��<.�IyTBhnn�X��z&qj]S��MR��4e$�K��n��
�,��
�Q���AE���E�߽+~)��'��q�Y���$kua`��#�G�Q`��>��s%�ـ=�}��\��dzc�R���˃�cJL�v���V�W��1�c�>ϓbJ�-�y�<P1EQ���X�m�Qc�䯙��b;vd��ʦ�� ,[�'��C`����D| s����)'�e�R���4���,>�g��`�u&�A����I�쑠Ȼ>M�rh���Z	��R�(������֏����\��w��C��J'���524�����.Ʀ�ϵy=4�1�+����[�u�kP���c=c�����\�I�����]�v����|��P���[�t�u�CNd�M��q��ȳ�>��E�H8�zPD