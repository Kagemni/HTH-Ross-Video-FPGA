��/  L�S���]��Ɗ�;�Y$ �aE�|g�}Tؒ_�%ǟe<$����.f;p���$Ǟ�U�_ 4:�n������ý+OSU/��{�֌xE,���pc5�A���ج�(�B�G�,�����5����:�rv֯�W�ֽ&9�����CH{����nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�UtK��^�)A��LTcmQ�d->m}oؠ�t�Tԉx�<�cB�f"��x��0��g�����x��z���5V��O���q�Վ���P��W�����c�^��� ��o��J�H��k�(|'K6j����3O��a�\�$����>Mu�	��d�������	���|�"�߁'D���[��^���ŋ�nb�����&k(�x����Ȭz���خ���8㞣_�w�)��j8�/QK���Ǒ���6|����ײ��
]�)����F�r��	T��Q� }Ӝ=?��c�@T��Ņy^����̙�ȑ� ������-�<n�''=Z1熁���j���h�QĮ��]����8�vT.WZ=�lg�[0����vm��t��s��K�ŏ����Yzp
�b8�{��dW ��Q�x7��ifp�m�<�X��8f,�	�Α�4ɞ6�W��.�j����.)1�Ô��I�N$����"�{/��Ke�t8U�M#�<���F^+)��Yn��^ƛ¬��E�[u���:	%{�``G��޹����d������Z��ü�b���yr����cڞ49Q�`-)�n��pI;G�?���/�O�%(d�I6�o���cz���oP�����9�-���(�u��
=kX<����Z����|�R�k�0�"�Pӷ5[4<�epN�~Tt$�~f��g��_5}yhL?!hH���@���Y�.�Z�lO#,b�A�{�-Q%te�s��2m��%��(x�C[��K��:�oP�[��u!���}r}E7�q.,HO�
1���_�l���dF�N�n��0g���V�s|�c2z�В�?�F��w�Mlx]w���	%�Z%,��$�Ƥ ޥ�@Ī��3k����<���%�ٳm��
5 Y}r�=Aќ�{�V�]���A�%�X��j�2��g��`ё�WR7%hJ��.�y���!�=�)>�6l��jQ���t�Pk+�kھ��t�s+u�=�M��T�utd5 e������V�+Xv�.2�Ѻ�Wa�����<Ģ��ƒ�#MWl!aP##�e���+͟�`�Q�t音K�����^�����Y��Ф�_A��N\	��}��}$�z�wR��;��k\�C�������r ���%i�D3/~���Ô",�Ox��4K �w:�_�v%�Z� ��G �ҥ��)�C����l����{�-���E�3=Y�z�7q�2���U�����G�Y��"�$�6����;y�n�e��.�]L����o��oWHНN;��b�! xHf��
����~��������"�D/ɍ�Ťճ�$��h��_"�9^������l���H��)H��=!Y�x���-��5E���4�Z�?n]z�K����c�SQ�G�Px�xcٯ�dzFV*�U�~���+���Q�a����5T�h�$�V�M�{�'�v �a{i����1�F�@��Q4#B��gm�ǹ��C���~���)̮7BH����K⮶հ�;Cɪ�)��:�_�G�����o�,9�EH�J����y��^T*�β�al'w�^�G��)mY�=^��E+`79��':�E���H鉎��ri1md�|�����{=9J>�Sg��X������$ZF�Z���o���(��T-��Dϵ#4$��W�y���)2B61�vj�6�Nm�9��_�~��`{Pʎ�=v�'���G�MQzeKC���T�qvb��Ī��y#�Ǣ�g�*�M��u���w�<	�x�v�����0��hO���b_)$�����vU��3�I9B���e�H�ԇ�=�7OY%��-=^��D\�سLkV�Ȫm���n�K6�|�]�nl֚ ���b�Hr�����H�i�0�I~u:Q�6סH�q;�j�|��Mh�����N�}Q���}ԉ�o�.5D���%$�H$E��˝�qz1��<���1An�ϓH�v��ʘ�%Y����H�T*q�������]��@ԩ�4�t{�»���8�𽱨jI!�kLG���T�o�'�o�����ą���.��V��瘬��t�X�@#�B{����ü�kp`�K�5\��>ɞR
�+��)"6B"����<t�ؼ�������%P#W��S+R�0s��`͌�<<���?��8��!��=3I����?�H�蔝����z���G�����*'�.�M���C,�QT����Z nG���8�a��}q�|�I�赽���/���`~�F��!�{Q������Į�@�LTY��aR	Q����$�z�.m����/����̛��$�P9V���o�d�J��������7zW �BE�^���|�nя`�Vj�)d\.�A�dF+�q�Ʊܣ�b��p�Y�"�u�!��?Ll��q��n��˯���O��DU���\�q��P�Ƞ�łrpx#��H�E �8���#�)�_N�(����[i-�C|�Y_�������������@��U}Z �*��yD@q�R�gJZ�}W�/����4�,�`�N�������G�����+��ww���7h;�);	V�LC��P��a&G�X�MӖ��htʊ7q=Uy�,ǉ���#�<z|4d�����Z�s�����_��U�%>�k%w|G&�ɟL�X-�3<kfe*����I�=�,�ڽ6P7漣D��J�0���$\
]��׽B;�)eS��dD4(�y҅F�W���!9������#bBs�V��^��1rN&���-�,>D4��3i!>ZF��M�ɵ�;J�P�w,_�(�h��i&�{����M�����!HdNtԺF��A���}����1��wٶ;�JR�Lۡ[v��A�rt��,w�}OQ��m�[ ����U2V����C1�Xa!_���a�*�"]>����':z���R`Q��Ñ�'�<��Z�pڈk*Ԑ�w������W��2Nig�S/�/�r�Ҹ����"������.��'�����4�$v:ф0�%djn0�5U����l�[�����j�8`&�b�����߃��dp���DUUP�1M���s�">���׀+�#Ψ�a���B�QF�:��}��̕q�{^9��K�+ܴ�$�����L*&�RŅ������A�	H9`$��S;��\hE��|gyN�;��:�������323dkʋ4*D�F������X�Cd)�O������CǤ���� }@b�eY���p-����LK]�1�</�� M���T>��x���q`��?����k�Jt�i����
Z��.�#~+��tr�֤��]���r�zrT���&_���}?]�&�J�Tw�=Z9���uY/Y�,��w3����6��]��D���_ܯ���X�e�X��)2h��צ�#��k���*^��fn�^��Uq���n�ܥ4�^�-�qH�X����s�<�
�Mۡ1AW���k�A�:�h5��}-�	��X:ՁM����@�bF������.&����.����'��;�*�զQD��!)�Ѳu�jY�i	�;�5�U?�
�}xn�VH ���E3d2B1�fu�tn .kЂ[�T9�b��[���z\��hX�I�y2�x>�fw����I>�Ç[�8r���	C���=��o`P_�Y��t-����H���<�y��h�"��W�SVĪhԡ�s�j��V�};̙�{ݴ����>k��@�ov��\�E��;��Η�O>��� 7�=h%�t�:�B��V_�%5{]���5����V��|Ae�7��xS� �����O��{��,`�ߗ�)�d�g��~���/.jpic������-�a`���D�E�Be�;8�^�*Ub�	o�:���͊B��G�1���m�j
�}K���m9ٴp�
@�f�M�����+�RR���%���	��\c��"�~�h��O?1(���N���R�Ǆb��\����H�������SY��I�;��_	�X�L�y��e��tg��g?��'�O�i[YQ����$ ]�H\���ȅS�/�4g�<4�׵�yKYX���O邤�/\k�\̾���y1G��X�-�+M���j`������Ϟ,W��]ca�X��Dm R���y%�^�N+�롕�r+��I�&u�|C��Y?"�b��f���J��J�����Hz��i��Fw4-ֈiS��S YBo�12��-z�������� w�AV���%����]*��e�No��|�:.5��Aj���LÞ�g+��L�s�#�$��H��z�+#2�1jޣvɳ	�Y��Bצm�B�� г�����o�۪~�����F�"��ZS>uk�@��n1ӭ��`y�A�h�7�v�鯮ˇ��"�l��:�����y�sR+LZ#&^q��FE�d���Z�T#^)���ŧg�*�Dqj8Z�U88��݃��eg�LwG�sۖk����^Β��%�+����]T�uf�TG���=�bEA��њ�rl�tG��8��0�`��p�-�!G�Q�U@���G�B��c#ߐ���.F���
V�}�(�
+B�+�%�e�<H>�]w�s����>��1�½�� �r]�j�u�kX��q�BM~`r�%g|�J	�VD������Y�e�h��I\u_&N��=E!%Rox�����ݽ���Ag3����) �H���Î��I�I�)n� XF��w��4cX���F.���