��/  ���>c��>}�r4��GL���wV0����8�^ϋ|7=b�C�T"�K~R�a�!Ǌɱ����S	"B�P騈��
�:��ڑ�J��^w��*R#��:�|�u���;���.�<0т�`~:/�RS���*;�X��1-g|a�ӷI$P"�����nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n����D3ӡ���p"�pM�x �GIc�W�	� ��S�w��Jƙ�����O�A|$a������69�nSd*yq��2��q��V�Qġ?ϥ�
MiS�v���$q>��b�P/�e��\�Q�T�)D)�W�:3g�V��[4���f�u~�Y��ڦb�B��e�XEh�h �b�m�U�"�Vf�
*T>P͛F��*��A#^��>���x��T[Oܸ���[�"����W�w����ޔu���2Z׋�{f����e�&W|�(
 >.�e���Yw	�q��m|�4e�'� �����l�����l��$F>���q��~��ul#
%x��HzlCFu�>F����}v��sz�Lf�V�:��IZzcT�(��+~%/�Ǟ+`�˅��a��k����QaAڋ� 	!��5p^��9zq�������IT�=��IF�<`1,�O#��R���Z��@#L�Kq{�|D�i�۟�����uM�i�l�L
i�8ٌ�D��na�E
'ݟ^�KEi||*���8L�Zۧ���v��4[3B�?iN��A|S�N��������v���Ru��=[�T��g�l6W/QJ�D޷8�
,�)��Œ��t}7�?�4`cs��Q���k�LP;���\ɉ3h2r��.�*L3EVg�
�Z��Jy&�T�����ۺ�o�P����׳��6�rW�T,џ�8%(�Y�>�$�PY$�ѭ����U�R�����A漊^bE�j�ԝ��]t1�I �^��=[*��P���(�����q!�t�������,D��:��EkLo�r;:lt4��_�}�ǐ�H�
,j�^j�V��Ά�܇5�C��=P�q�L!��EO�P�bh�ó*%{�ء�Ÿ�	�LV�F r^�Z��\�A��ҝ�������+,ek����jM���U��*�\�˙��tE��~�Y4���5�(e0fg,%b�����r$���Et�24C�J�%��B ��Rj
0ւ�߸ ά\�)���=>Q#d�B��
��:�*q�N׹�6�S�'KWRCZ�#�$�(��[��X������a����:=�G�?���JK/�tY�`  g�V��R �0^�����9�h3z�Y��	c���#&�.Lӷ�'g8jQ+�B�,�W�EA��$�?b���"t{����I&�죘(��p0Ü���V�� �S��-/�Ⲇ	:�B9
�ם�X<��d��l������G!a��^h|�Ǚi��C5p
�'Zd���8�$�I�R��%�Y�.o��x�루����4c�u�ϥ��A|�=�{X$������'��y9أ� �}��a{,���(�����O�P��4��r��n��.���������|���Ig��^R�xc�H�@�Ss���Un��G<��@���-Q���?�L���[�3��:uɗ�� *�Mȱ3Ͱ�������[�t�g/�h�R3���҇���|�C͡�爌t��M$/ڮS "���,eq���$Q�lp�/������;��/�7��}�F��8�Y6���6�E����v		�G�?�KzU�谬<�����h�Xݏ,�C���ټ��zdsk�ПO���9wGm.�ʭ��l�EZV|E�>�Q`\�j�-��{���[�ٵqh�{A��d @o�d�@IymNƘ�M=#\P�7��0ؽ��2��������a�iލ؎W�Ru����f���&�:4d>���IZ�B��PgVz�xn�dx�s�v^+1�6�X}�ɵͱ�7P���"�B�ǰZ.�pf���gHg��z��)�r�<�>Q��iܗ{br�QE"���e�GqBt;R���@� ��� �W��ג�Qm��M��~���QMT*����I��j� ����|d<{�U��%�zZ�d&���5�$�%s7#��ܨ�$t�p�ŀ� '�oS�IVT�_�n�d���7"u�o��	���bo0m?WϷ�ɵ��N��<��ɥ'���D�������0)yz��O6�_��f�7&A2�}�B��Bw]�nќ�~�A���m����D��`DO]#�\�4(�< �E���߸~�����K���a����I��q����qĊ�$����N�@�n����]��b5�^2_L:���T��H
,7�%�"�Si���G�o��st�_v�P\q��x��vD���_"�؁������E��r}�&V{?*S�#(d�ԏ����+�E�p;��}83jya�@r�a��L���}�͟o���m��Aل� *��N3�u���L��G�e�}-\M��4[6�&�Z��1�� r 킮�B���;��m/eG
6��������§���c��j�����3l{�RWg�ߔ�������)�y���R�4G��y*]��|�K��LPbH:K�[�\�y�Oϳ1�$��� fX�Y���$K��q���S�[e־�M�{�G`�,�=,�|\���p�D�g�0�R�B	]�
�V=��PY�&��C�I�t�fN|�/�Të��F������S�<;�]�R����o���h<"������� ��5)i��|���fa�Ǡ�<u�)���F�	U�DL������A�'�-OzO>R�{L	���PEN����+՞-ֱ�n�p,��d���c/��{v�ܟ�.RpI�-]�d@uB���)gO�Y��Sӌ��CS��h$���[���˻�y4��л����&��z �����I���3�q���ß��0`��<ߣ������׌� �Q�<Cg�'����g�]
���s5G��mg�{t �YV^\&[�*��,���[U>aLvu��HO�H�?~�aB�}�쓹X�a��'�C[�u�Rd("���,�����(��r��<������>A����(-��Е:x��T��y0���ʰ6��VSE�|����7Յ��L>X+0�%�5Tʘ{�G��*��]�����m�ݵ�F#,"r�����-`�u�#CG�aW���>�󺟭.HQ�T�d�?
�r�Z�3_X�M?��N�ڲ�C҄��_%[s470�I9i]��=%�#F��Nb�'dj�˷�%���`x�A�׸"�����}TV)��Ejq��]*Q"�IhϞ/&�=ߤi�� ���oɔ!:M�O�V�T�d���r�+v���`�Q��U����K����հ���F���a�NZ�*���V|��)ު$Mhb��|��� �d�����ȍ�/�h(����/�^�W8�4T�B�=�ˎMZ(\_Q� �L�E/D�E�enR3��Ώ(s���F|����|��z^1�{#@$L�i�֘�m�z<�\B�<��/s=�̬��ü>c����9�U9���(6�BQ���S�L��b�'3�%<��}��V��F��V�'
Y��l4� �I��pSJ�$F1c����
��<�P{�2vrS�]E���o÷��KV�B:4K-�G�y?��֐�|W"��r�n�ނ����q5��!���H��J�G\%ޤ�<v�R>���s���%���-ՠ�U�Z[����NA�z��ղ{�qЋ�9d��uG��e���;d��ڧX�����cc��e6��F]g�vƥ�Z�f�I3I�-�����C���+z0�MU�� Q"X�Ӊ�c������?C�BI"�7�5�B�Y[��4TQ� 3�i���RG�M�8q�-��l�k�,�b�8�\1f��e�JS�,xr�/��=��o>#6w`�_H�	�w��2���ԾH�&AF�gy����x�Q�$i��P�h|��	��2d�5/[C�n\C5Z8�h��sLd˳R�a��ߕ�����ȿiDC�"�2�R��˰ԩ��P`"�ٕ�3D���qM�7hA��}p#�5���Q��eŌL莯���ǡ�� D]V`02��L.[�s�-�զ�'���Q�k�ghR{�i�}&�˕����B�M�_^�L���寧3�jj�|�%��w�}�I6�"����s�zeޭP����=���Z�p���w��^�,����|�8�o+�/����[�vM����Ε��n'��́t��E���D���$|���a��x���L��Ɖsg#�9�0;�K�]A�/��$	@WVhM	>B� pƉUn��R �C(aQ�ǀ#U&\jo_��2A/�,k��&@&-"0X��c�\��yX����8JY������]=�"�`5t;��:R:�.������ȫ�Gכ�6�ڶΰ��F5�n�8>��AH����{pe�f�P�,�9x�i;���n��2�a���������Ul�c9�fi�� �_��{�B٣��F�$>k��L ���"b��G��ǳ�>�{��f!�xsbOu�A��3����6���'E.�rВ!��7¤S�J.B'v��w�K���vF�{?$:�\ ��nEys�{���_ˈq�8')��:d%�P����O�W��k�jS�p�}-k'����"�@��j�l�Rn��Oj'�b]Dz�`�d�G(רء����>��M�]kY�,%�IU�H�a��.S�r_|G�L�RONv��H�W�5+P�s&�q���,b`�OH��͋h���d'QW�mJ6�'�B!0Gc��		�*�7��E/W�7ӽ���}�(Rݜ{YFO���4~�ٗ��X�	P���ZZ��+mؾg��ip%�(���5��Rf:V���A��~'ˇ�9k�3<��-C/mz� HS�osR�2EM"c�*��)֬�����6w�,K��Z��R0OT����wU�����}46z�B߮��_������ox��&=k�Q3��+�-�Ю<&��_�Ɛ*�fǈ������k����ڽ]-�>|@��`�������e&���F�[�w�E��-�fB�)�'C�k�f3�ϟP1������q5��X`��W��+饨��"�q�.��y�u/�e���H�x�2��ݽV�*�~�F��I��wn����fۼ&}\'*7����#�S@0�mZv�"Q�)/��*!9	,���$qLd �����m�65���xӯ:!�z8 �>+	 �BQ9m03\"�|<��t	,X/��94E��Ў�QD�7��27�L-aC7���3�h��]�ڣ�*�k�X�8��x�aqx)��^.�i�>$e��)c֝t8/y��>��½}��%
(��!�g؋�3I��2�<_`d��7%��c ��v6벴�V^aʀ8���(��:��N�B�Cm�"�Yi١�� �?��O��46�*����c.^u�3������/G���A��eA&�ѵ�Xn����h ��KP<�bӸ�j�+��s��ք�F��uq,=���`�����6�-h�3� =�_��޵<�-(~�n��*�V�iNVg��0���$�J����
.���oS3��R8�0���YP($.�՗Ձ�P+)�`��k:0���O�`��{���D6�e��*�c��լI#�qWYG<?E�։�:�~���+�.U������F����Ț�p6�D�ȩK��	���AZ�0�9�
���=�[ӟy9TrR�Z��ux��.u	)x�`� �x����u[#�C(�� F��Hp����8�j����ĐO�"9�l��el��w��-�K�NJ�%h킺a{���1|vn=����\��V��'��VEڱͦEx�o��wz��_�Q>�c�'ښ�N|���v4ѨT�֠��y�U'��|��0�v�$�dYh����ܦ�T�N��4��dJ�{���n(���,D��㤗���wy~�R��f�I�e�B�[�4�)ߖ���[ض�
��a���� ���i�{�Q��t�b�z]wA�uo���8u��hߖnC�_�#.�~R�F��*na� c���ɕ,����zBS���X��9+��6�K�
?��Lp���	NEB��y9���A�+2�+��ڧ���� n��Ǖ��p�ۘ���Q�����R0����sHޥ��k�jٛУy���ذ�AtO�7���i-��z��j��6��^���|���N�v\�:'�͟�ڢG����~"� �ěG�r^�'��c�oy�i�%W����0��-K�B�8y�R܀lq�(Tݚ�fv (}r�;(m�B��^"Y��O�왨+��좴�>��$��dw/��E�Ì�7��4�ۋ[T���[~��B�1�J�*왑���J%��es�¤&�t��o���C��$Ԩޯz�Y��U����58�:5O���znHS�f��t�DE�K�ro�a��~�:\i��iO���?�'�Ǚ�k��$)��P^�i�>,r)#8�1H���ɑ!mA_�H�܊�&�5����@#p��c�R���L	�$�]5��rv���Q��j�&��˽<��+us��V-�z[wQ��&P&����%�n%g��i+ڦj<c�C�%��ߎ�gq��1��h{�U��2ytU�_�<�Sg��3���ܾ%s8�}P�����836g����"�|L*�k����K2�ٽ�̙���k3ai���h9�*�O�V����T�8BHp�ͩ�c^2C�^���&u�s�l�ط��)�)e�t�i���kQ�|���������҇��U�@$[�Cm��A���8h���-YAH\cM�ɍ�W�0rK\��:����B��O@��0�gP6b�Y����Մiׅ�,�v4��^Z��g�%'��R��߹�[U�����G�W��Q�$�"�I���,����@��L7�x	`i�U�M>-^O����,��������FH�I��$�"�LK;̑�v� j����A�2wv����c"o��j9��?�L��b&�d��j��HϏ�����?�A��ZiN:��vj��0��o�F�2�����qk�WC�?��L%��,P���rӵ�H¶�
�ɘ��	<,�'B^D��x�Wˣ@&����a�[$&{�F_�?_��w�3<�ھ|��>�E�������Z�g5($��.ܻ$�z��>B�8�t3M ďB�<�g�PZٍJ#�J��|Ő�d���E^~��p��uP|�+m��4�R� � �O _C������΃C[����p���LǉI{;��<�H����}2�I�N����Y�г�Gu�P+z�_òz�����nD	g+Ά�@K_oj���;��Ya�}��
ni'�'�����:�ʛ奟���jIȬ���Ĳ��{�Ͽs��!�P��a*#��բ+�' ��o�kns����*�c�,KgA��87=�"���dJ�o2�e�g�}_�l��Ѡ��u=&Oׁ	e|qAj�2��}� D��+�_m���>=0� �43%&n�ފ��2�h4�T��E}�ƨk�6m�]AMv�Q������i`�)D�U�l<�;+U��h��@����w�ҵ_�D|�F�h:��������c��N��g��4OEŀ��&, 
@�ߨw,�0�|�B���Kя�u��
퓡��=��K�R
�`�!e��$��D�:�9�@-N��s'8P�1�"Q���!S/�&���Ik�\z�О��
�߆N��Z�]pG��e�
��� ̓OG7���:Ml?�}Ѹ��Bfb2�f�ȫ����E�r�i�DJ���k�J����fk����"]#/���'�eȑ���bK0�Pձ�Z���M�Յ�4PKٚQ�Ȧ�뫮]�*S�?� Y�
���3?%���A�G��3�Z���\}���s�M�.�Z';R�Sc�"�i��Fҹʷ*6�Y>���-�ݷ��K;���g/�Cw�ni�*�7u�T���
�"�l ���D@ސ��(_��3I!��u_k�A6o�5�<g��*<{+,�'���:v���wkp{��(",+���G%��;r�Gwsz$"��7�h�]wd�����9m?�0�٭8��Ga�MXl(:�d�z;�LL��'��O���;����_W��j�I�Nu�� ɑ��k۱-������H��'0���u
*]N�3=#�xf��3���a���]��:��H_��AȊ<`��~vT+�9�`�͋5F�`�[bT
��h����1ReN��08��,A^�i �]=�������!s|���������$�
�I�@�֗:��V�����z)^"G�0n�\�~Z�iҔ�"��jof7�q�CA$�w�(��L�$���I��`9"��t�*�1#�Q�	���ԕ�9H���8ʼM8�+_yF����H�5<jf�{cBm�eѣSnR)�&+]��V����!%�ݸ�<��]BP��i_u	ʇ��
��W��t��6�@y��Mz���m� @�Q�Ʌ��煋��a��o�H����[�z�x
ryǺd�si>� 9I9Y( ���5?���:�|n��L#�U�(��å�S�b��r�_�ۤ�eY'y���c�K�d�=ޜ�U�|�9��FT���7:D�H�옷RP�*!���	� ~H� �ECl��{�����}�lso���o�$c�5W��@r�/msǖ��yh���Q����Xߓ#�yH�;<d%�oB���h;Ff��1����ôT)/�Z�@A��_18r�@��5��d|����^ωl�@:΂���wZUH��4�����fz=����ݮ��L8(,b�R������C_ф��i��^��8~�����qNoQ�v��$���~+�F��jT��їi���RdW���N#
Zf2ret<ӖTfS�0\�Ox�,G��� !���|'�T��q�;�a�� �����n��;=.��������T;s�>-*KшEo�uR� 0;��?F�-,���@\��O��&���&�B��o!�̬��mP���-*��Ż�uA�+v8v�w���S7���g�ऑIh�A��
�~ ���K��h��&l�Z�W�:!�81�I��ò*���^��2zцQ�As������J�'������a°���O	Ҿ*O맬����|�Z�p�ŧkMt����J�I-l��o��K��W�J�57�rP8���s���1�:\���"H�	2����p�
 �!h���_�W@��gt2c���FtԖy���3턱��נ���Ы�`�;݇��`���XO��ᦔ���
�|ŨÏ��z�Sx��L���di'�� A�N�y���Gg#��-4D�i�QpZy�-�wYh^_
�)����$`��w� /N��V�a�aԥ���ڱLE^샙ڸA�&\�qh_�����=8��4;*�ƬwSjUqN���q��bu;1@�]%')H�M���PPh�:>sӃ6��#��`0 "�*��)��U��w+�5���G�~�a�/*\���{5І�����=PM�<��&A��ġ �F5{��.p�P�j���R/qs��r�Q���=:��5��.b��b��p�uB
��.6��z>c�ma���3�v�]��H�i�S��.�m	W}�}��Xb�������	�m�	G"�J�2���@��� �8�?��l���k$�!T�"9_�6�B�?�ڸ7��:�9hq"�U�J'!?;��%���ⅷ�