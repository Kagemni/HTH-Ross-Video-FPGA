��/  Gɭik�ﶫ%ū�Xh)Y���:��u�$�~ zf������+@�CT7��R�a�J/��Ώ���CF ��:�`�5�-~=_�*Fowx���(�]Mcx�D��Rt \kg��T�����?'�Um.�� �F��M�ǈi����rF����U�)�� ��+'��a+��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n��:>7ߎ��Ғa��H�Ɯyї^sXz�1>l��^OɧF�e\p��.�Բ�O�mVZY�5F�G�����"� z�mLb��ă� b��o�*|��>�kOLt��z�(iR}z���עg��=��\���R:�ny0�;�J��ߧw6�w��e��`|�4�~� �����?Y3�A�D�λU{RMul�p����\k��Z��핼󕋵\��y���cm�q@&���I��Y9� T�P*X��͜I�KBp�����8z�6���A������~Љ�w	 L¶����������2�_j�!��e����+l�X�I�ɫb~�r�M=��0O P�����X�1{�����6ad@c1ˋA��M~�̘2p�i�?�b��?솜�}��WV�G��Q��}e��'��9f٬ή�X�"��j��閖,��Ձi�ƚJP"P��	!˿����v��^ѿ��6��ٴڡ�OzM�>tbe���xd=&ԑ)&?G=���w�:��F�s YA��J��a�"և����)���I�h�^��19�ܴW���7�ۣY7�!��	xJaFk��	2���dGv��S��
�!��D���Kb�d�/bqe����=�)��M�<��V��OX�Qi��3��Sv��a�@���H���o�9%�I,��y�m,B�T �xH.�|������'��%�赊�|A�����6A�Eăn��Ѵ��a6�
 �'���54u�?$��7�� �SY���j��ݨ����c�K���3��ͽ�::�e@������Q@.��B�[��֋��$���ҳ�:"�Y1�:�Eb#f�"��:@�R��\p�/>7�����[[�+�$"j"���~R���bz�9,cGv��2�
T�/�4�Y�?��Mࡊii���u��1�ު��&�q�����q�pj+J�K���>8Խ/x�a[�s]Q�Լ�k����Z�B�f�1�0%#گ����n�R�1L'��Z�O�UD
� �w��GR�"�/w�߈$0쨆{ ��p<_���e_u����e��m>��/k)�y�\|��U�{Uu�C�_�OC���*�B�劎T]�6�ڊ��<�U�6�<���R�*u':Bh�l@�?��Җ0r���(� AZ�Q�%�fޅ��@.���x'M�!��nE�ȥ���]񌊝+�3�	�n��Ä�
I�Z��yʤ_l-�x���Xa��
��ڞ�؀�{���MB�OP�M���L�E^���Xwy��O� -��!L΋G\f�T��W�� ��n/;8�l@�uƔ��7֒�u~LzVϞ*��i�q�o` �Գa��$mt=�$N�����@�?��s�	(j�|�AY;�l��O�'���j�zL��p��w�x��r@QJ�ch��I �K�|��w���m��(u�b�<�=�e@����!�����٪glÐ��2Y�8�!b64���rJ���$���B��Ʈ��h�]���6 @�o��Y���������A��������Ȝ�4� �]� )>��� ��&	Qq����Q8:>�k�=;:��MC����.0����a �0䨅�(T�?=v�����i�X[>�h�<k��S��o���B�B=�F�K��_�VJ�}�m���-��}�[O&%n���Pz�kf��FwwOP�	y>0[v������,ĕ3pmdz�mr���=�tʯ�rϩQ�D��Ke.�T�a(:�Fw@���0g���1�����Q��a��b��r��u ko�Т_�o�Ijb~�܊�P}�(-K�����G�Zl����޴?��\�̖��2�^!�z��Y��9���?�S=�;��hV�3��9����]��nw��)�.�t��=�t���X.p�G�.0[������ Z���
c�h
��a��|�G�S;mw�gڑ���&���N\QO�+����;���P��j$p�KK�&�U�OD(mY!�D��t�)���2��F&�w�S�IىG��DH��OcT`���D5����±v]8]�,	Ҿ��{����x�RK8G� o%=h2�ks>���ItŴ�zZ���$P���y��ŀ<^����(����o�)��D�1]AjY�m�Q��Ӳ������Y��?���d�`�;�?WV�C����f��.U�p���-��sՊ�I�ƄjH�S�eE�~�7��b%=��s0��y;�Fuh*�},,�PcH �>B��+s��q�n��KAF������<�96t�rT#��4u��F�Q��X
s��1�,�(�R���x�u}�'jaYt�tĠ1d����3��d篠m}F���#�?��yq��f_$�'���V����Br5��0�GVix��h�q����W(�wMW�~w�ws��ȤV�����$����h��
�����Rm��ϣ1�V��'��7��rK�\�.Ib� q8^��\1�.���a9��b���P^�yeQ}���.�ѣcB{�-�u�I�w�a��O1k�}DɿN�!\N�����[ծ��E�6�܂�0q�U�ԉ��?B!(�Bee�NS l�5�~Z]ŬӇ�_�@� ;��u�\�)pi�y��f5�!|�_�I��s-'�i����(J1�F�&^����5Cߣ���->=�ut[2��#1��~���L�N[��t�trWL�(n�ҹ�
�I�#6�s�.���iġ�67��G[!�b�T�7ݭ�	2k8g�[P0a�"$'��1���5e,���#���Em��ٍ��{"gaN�۵1u���QH�߷�'O�❙0w���Ш��-XG�$|�+m�0�������z1ޖ?G�S��t�,?T�K�,s����%�Ʉ�u��?ӓn�t��GR����A]��<zu�����q蚸Q;��H�`�(�N����� ���L�<B����@�1��f9{(�������co6] M�	t�.G�-�ʖ4���P��Ƽ��[ȕ-�Ao����pa�uAep�bv���~&��u}\J�[ۀ���C\�h*�P�d��YM�C�!.��c/]���ԿW9b���cq=L�vW��Usۿ���ʗ81�S@2�B7ګ�T$��0�3�L�p��,iPsz.�34�~/4�`��\nwb�^nb�B�;������x�ݟj�u�d�0��gW<�����Ԏ�&#��w��绐�D'P�/Fz��u������v�>�����o�A�,!�j�`�_e�c̟oL���e3�eH���:O�	H��.��
��ę�Q���ff�Rwm�x�.�J�Z���Zo�~��;�}ֆ����&�O�4
�������LJ�3�@[�'?OM9gs	ۛU��%m��n�GZs��}9�+�̾����'�}���rFa�EE��E/	�a��8u��{(rd��>�q55���b&R7��:��V�	��Kk�V��$��{ʕ^�I�B�P�M��!H��k�v8�����E��V������K\�<�o�b�'j>}��>ϵ�V�K+o�0Q��?����Qw�B���+L|�� �$� g`��Eij)�E5��0AX2����/����HZs����]V5�ͤ�
�:q���Q�%���b;w墍^pT{�%A��'�IC�i9���sO)�����=/����Vl@�>�U�i
a�q��[�p�<�;YOYT]U&��ז/_X�R ����<7�m^�`F&��j�Ȩ�fU-�F37�z2m����J�G�� ����n�n����
L����\]� �@��9,���m?�kP����s#��CMd�9
²|�i�L��K223�i����E �@5y=�p\��d��5P-�wU$�U�8���n����P��m��е��k��]o^���!�7[L9�9����u<,0W��?��c�}2h�MZ���0�i瑯�¹�������4����XQ�쪮(f٘G[tͷE�nI-�D��K�͓��~ueb2�k�V)kP/ТNɬo�]=T`�X2�5��ܽ�T0�F%�<,�����3f��
�CN,�Ъ����ḫ�M�{
s����Ε�u���n����ߒ_��]uQ�[SLM�F�W�:Q�{Ƙ���?'�Iَc�<c�����ѭ֠@��� T��ʸ�(kߤ��.���Yv�t���Jtǻ�J��|�=�c�wBN�fBWG�.cdS:�xY����I�Q񉩳�) EA�j�ђ?�W����f�  Զ���,��4rj���iS����ڋz���u6$�"��/������Y��1\��B��Cm+�=2�D���1�5kl~�Cc�tB��h�v��J^���(����_aN���B�;sw�BX�51�NAz��-�4:�Э�'MCj�m��ps�P��7֩�k���yV�(�t�;s��֐�Fd����a^�U{yya���z��&\�i�`Y�0>�l�e�Ow{�<to�;�W�wk�6i$����<��
	Av1�(��Z�����䷹���
����=��<�����M�O���!'�(LM��O��`Y���׊}ՠ���Rq��b��N�nU�S]�h1wZ�X�F��)�ʌ��5$r�|��F�����y൚wc�*6K)m?�Yo������-��FFgǕ'����}'��cq�}��+�̨���z�ݹ�3dm3k�ݧ]��,	�1��of?���'�)K_�:��{xE�aT��=��1!���l"�����G'*U��݆a��[� �=T��Q+��Օ)����a'5��z��cU��m�Ơ�\��I��R/�Y̣�c7,O{���U<�k@O��x\��N�E=�
��Ԡ��PuC7#���,s@��D��S���<�G�p���8���C��|$�*T+�\BYd���vB�9ʣ��f�@~獥f0���N����W��v���uz׵5�j��MD^귺�z[f@��p�	����;$�y���G��Yr4d:��8��H]��F��}� ��Vo�p"��'���bEz2�T>bIW,]a���^����aA�~36E	��9�����߉��ED+����N ����M��ҿH�Z����ZB�8h�]�]�7=���?>�eέg��X�	�"�C=�W0��� ~YM���N�͐'��yl�J�ܜ�Ҷ挘Nu#^B��l9 }����{��=�p� �d��G��W�}Ҧ�U��G9�u��g���]@Rg?�&nC�Ė<T5��N|�k ��@��Y�:�O�2����z�z�gFv��`n9Ht�t�'��="�a��+�9\eEt�H��t]�4H�xUM!+hn7_R��5�.S|w28�����f���ZҔ���r�UNc��Z�n��X2�(K<X�`ɪ���&S�`���/����bf�Ofʮ&}w!�;��#k�]�x1�5�HM�^�*�h��i���J9z�+�
[Fil���Pm�Ԓ�-����;�����ײ
\����|Gjx�O�wO�ҽ�`	9����J����pG��(U�F��l�JƝ�_W{|���Q����_1Њ�昔���y,���X$�W��l�Ru\?�ܧ�1�ћ=���쌡��-�$�)�{���q���ӸoC��5�K˴��R֜DL��|؛���&��0�B}�ö���i�0��EL�iI!�X�{bv	�^/�׽�o�+�g/�p�}/I���yyCsn��&6Ԟ��)E]�`E��D�4����>"���N�	%nVi�~:�%v���XXOB/�<��0<�4��}�LPI�Q�WF�eRk��/�/p�,t�Y�q�~����7�2e_�΃Q.bLVC����D�e������vvꀝ�h$��
�/�vD��	~QB�`��m���y��R���^�3c���
h�k�)I���?wM�f
���1�(t=e�<�����o��c�2��w�-��q�,�g��Ղ������i�m{A��"T���^���E{-�Ĺ����g*E��r�0�56H~��/p�4]��T�}Y:��!*¤ʐ���-�ktlI>�rҸ�WI���9����/I�0p����פ�T�$?�����Su�TD�aE�j��0������,O?�fƀg�������T����u#�ˢC��x��P}P��Y[,��Rd�*�|�Ğ0�Y�ˉʩSl��N<����(/Kh�����jʅ�mO�Q��� �Ǐz#�C�E4�!wTB�^8
R�P���Ț�d�(>Q���-H�,�R:��N�h����X�W,t9�O��H��Q��;V��t(Y�o�����WT�������U	���S<8�ׄ���:TnٺO���N#��
'
�z�??����A�^��Z�r?�%��A��ҡ�)ɹ���=�'��aa�Zϖ0�`��5 �����aXd�p�"��4>K����{!�d�:K6	s�{��߷2��q��Eε0ǧ�������4aնbٞ���p�`��p�@$X/*��ΏJ8 �R���ҍ�@,��-e�~�Tab�%�7R�@�ͳz���έU�F�㢻�[��<�\���������X��sQYQ�����q)�Ĩ)V�����H�e���ߐ�'^D�<u_�p:�z�:��=�*gS�{�"Ϥ��l���:�t�ЎX�d7����#�-J6��hH+l+���h�>��̻Ox�[�����=�����;[���P�|�]�kI2�K�ϛ9�'����п�v�����|yNU��=��7g���nN�hiM�0[�0Kh�| B�,��i�ȻR�+����ސ�}0��&��Aav"��q.��a���m��<Fa�%0�MH�>V�~4��/�,B��q��Ɖe�y
gV� m��G�=���0f@��yڤ..T�H�xDgXAq�̯Ų �[�v���I����ט�*��j�f�Y������cc�͠Z�ؿ(�S[<����ÑƗX���v�>ͥA���ki�.�6�����Z��8bmRհ!�W�j3s��E�R�xܰw��R�4lգioݰ��2�
c'�@��
=� ������N�+J�qo���,%� ��:�i�+{y;��d����A�H�E�S
���M�Nڀ�n	ڐ���h@�=v��B�DΜ��*5�f�<������߾�
|%X+�N��r���s'ԣ�h�w��H���&���[�����\��MX��Tj+<�(
"���{��������Q��-�Zq[�>���XJ�RV�$���*��ᅸo|��G���F&�a�3�	�2�q�nR�,^7T��O��T�ΘDÿ�`�}��#��Q�?�VHN����Vo�MQ���Y���؜�
�L� ���LoD+��R�q��E��#�J bC�G�d���������[ �����sMb%�R�2bkM�6W�y>�t_� V�r�;�'-��wB+�[˙��hؑVWk��杜��8n��(��]��^�y`u�I[Ѩ�����O5���'�ȶ�ܞHM��������	�%$��6�f�"��<�%��.s^&��[Yz��=�����"��ԻB�Mz�z��v�A���y�c'�{��~�R��<�Z�H=��1 �c%�G���<�F�����s�X��_ҚH����0u�����7�%H�0���%�z�A�}�_�(l���=�!C'��ſ^��m:��u�AI������/k0�f7�-!��%q�b���~��0q��P|̓�Fōg������f]ɐ$��4Z��V����c̹�;��{ܣ�14��H+�)}k�J0EK�lI�`��NN�Rd�e,��y�đ�d�B���7�[�7�����a_���tr(���Ok�6��O�J�AUd�}���[��s���܇'Z�9O�D�a�;oĪ<?Z�z�
kcs���D������et	8|��\��H w)�1�WМ]�� �WCj9@M����ք{/n�MM�#ʛ���7���.	�y	�9�͕��q�)4�bWYX=���Y_�dq[�3q3�9ڏJ�SzN�1�w/|��ߖaF��F\���	��9yk�~�r�{J�0��v?~J�ؔ���9�|p��c�����ݪA��)�ME7�H�ݓ�eNʘdp�1������뜌2��'_���w����D �S����2e�Yj_B�u �p�s�w+`�z$=�$�oĄ�o$|_�