��/  �^���H��Uh���4Υvi�@����m{Y��t���mR�לx^E1l���8��ꭠ�w��`�����ޡ�)�f�c��v+��'�WId�U�LUz��sba�!/t�7�"�>hW�g�{ i�`�"�A��^�4��%K��m�:�YU�9R�T��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�nG�v4�iZ���ÔgVwC/�N�T�_�;B���vQ����B�J���/�~�V�Iڪg���/&�r�r��I���NB-=�����Dei���f�m��_��>g�d�֯�ok]��6�SƄ nо�jN��X)��U򀵌���l�ƦJ�@r �$�T*��ݼ����l5j�5"�$	�3[���sX@��9�L��v �O
;H��4&-��j6��VzR>6�^;BwO5֑�rG�A��`���G��O�	-������*$�:��ԣq�pѐ����~��Tt|c&U�>��d���Z(�J�a�v�C���2���GR�C����ko��d/᎟E�k(!>�T�@�����~���s|f��K�Q&3b��]�9�K����RZ<8[�s�dHo�E:P�M��A6E�xz g:�&���W�X���^�U���6����4:S_�z|4�\�aS�dΟT<Xe��G1�,�f)����PcGo�n-SL�B�Rt�ߍ�J7�w0'4�P��� "7���ڃ�o��_�N�;M�n��3���Z���hL�<H/�f���_g���s1X��B\���K���s�H$��Ө{�Լ�|\����<����qe�Hd$��_��u�>Ǳ�>�NL��O4������0��0"#��Řt����Y7�7��\#��)1���M����WQ����&�	����$��� ��B��Š��gB1��H)����l�j��g EG�V�����Q�Alq��q�H|_�vJ�
�p*1��0FF�%*�c��7�r^��<]1gvw��:F��Ȧ����4�KMYVU�>�Lk:s5�+�n<xT�R�J��}f������bp25S��W'1���Au�(��j?��ե��4��V��\�#����6��� �n�w�SN&}"����������u������o��$zKR(��BM�n��5�5��Z�f�OјC�K�f���FQ'f��(��9�F#�HEϿ`>�9f�U���n���x]�W�����
{*U���(�:��7m�@t�L�֣�P#��?kBI%*-r�q�(�5�F��U������AǕ�����.OL�\�A�~+ϑ|.Z�(v��̿Y�r�����c���i�|j�Ah�6��ZqXWq'�K��,p��/E�`�ͬ#rT?��Cp�y�3&H:Oީ�j��b׋�e�uT�5��Xz���
KgI���x�
��:���k4�aV��G5���V�6��E�F�p�4c�b�4ߖ
�����ӻt�w}�f�|*-�y)�=ŬD8��
���T�2�[��5�A\�N3�XUj��
�,y�80^_��Հ�7P�f8ӡ��@��b~Hg�߆ $'P��(�/¡67�~���sH�/' qGL�O:��}�18`p�D5�uXi˥��us1��[8F��/��@uQD����:y���Z�_:���Y���e
f��>��G�����}��M������3r�+-�>���� E�Z�S���W��덭^r�o�z5r-F �V&�3�R��EYw�^���$��t[|�`;��=;�d��c��WI��8�@�gl"v$�H໊i���oP}oD�x��hW[�=_5T��U�\��u�{���8���\lK��l3�/;�q��vi�
LJ��9����������A;-��O/�P���t�n���0y��OhN�lq�N��$0�(ן`��<��c�?�[8|��ǓWBbfOz��¼��F���X�őj[!1��ʽ�C流�>γb�Z�o��x�`n�{�1$7�MOj���, '-���0��܏lQ��n�ZUI�����:���x?-퀫)`91�?��B��!�?5'o.��0$gx>z�� �}�1z�N-��1��i���*��;���>ȉf�	��Nf��R�1�i�b��V��`="3U��WΚ~b)��&�S}�LV4�R��J��tTOyU��}����bV�0}aG4�7�t�'���? d��&��"gbft?��Ͼ�-�������U/��e�����6ΟJ��7��t��N]�(�ȇ&��_�D���]��D�~��h�l��)�aK��.�yi}z`7�����$_��y�<��)����\���{3	g��ρKb[Z�I���z�:�~N��)�gL}��_����=��Ff��WL��N�^��8�'�\�pX��t��b�BF��u�B
p$��<��r�4�0 %���3?t�&�QEںԭ�%�p5u�4jm��Oz�z�j7��`}_?��&�q�cuC�0��H�T"�d��B�ׯ�{(��S%WNҸ2Sf���,g�{������ɍ����	V��0��e8,WoC������l��t�zr���Qᄿc�2ͻ����N���(�I��K��$0N� ����i�$v���8�w]�j;X'���ސ7z�S����Ԃ3�¤�Q%���r-%ڋ�յ����r5-3�i��k���s��W@��k��b������'K���b�2��ݎ�3�	�s�ZL�?[P!�Ʒ�~����13t�lԥ#��r�b`t��h1��<.K�K�%�F��QCP�!<�ꘋ�)s&K��}%Ɇf F��L�S��NJ�'M5�� �l FX�+�o���l�Oq�X��|�ʋ]Xy
D1\Gp?M:;�W!��i��d�o���NU�M%���S�*duT��Ο�Ĳiz 10�_�X�����4�F���nB�	E���XSO���)�1�z���1�N�
�bGW|�TZw�����!����JF��)`D})�
,��,~E�z0>B����n�u�ty��i#�ܯ�S4%�c������_����g�v$��J:�]@>24呮��~8��^��XӾN���}٪Xt�9K�U&�s%pm�r����k��T[?��̎���j�6��Չ�m��s������θ i�@�f0�s�Du�_nVϯ�\���~5L�`�}��Τ-Cg�/+���� ャ	�<�.�N�Lc�ru˵���c� i)��N��O�4Ҿx��ۧ�0}��_7���됊�k��@��qx�S'g�)�ɑ6�.�PŁ�QhԬ�`xO*(8�1l�Q�^'�`cL��B��NZ���ߒ�EM<�8<��F�yD�3�v�G�Ե�jw$�|��On���PE��U��4��"_�|��b�)�+P>�Qf̆���MJ�PU�GB���US�Њ���]�?���d�������,"�� U�As��K�4u�lt��}_��#��D 4���i�ohʹf��%M%���+iw�6��ǲ���Q8�:"ۿ9�Q��aO#�±�y��%���Ǳ.���3<G��OI����M�/�i��T�biz4�2���Y�]�^ǝ5W�6�P|3�N_�Q��z�r���l��2?����0oiD�Y���j��=�Mr$a������\��B��@W]AFF�6��>Y�3�ᏼ�l�q!��o|V&�<�.�%�5�	��*׈"}I2������]���D*�Ǘ��2�؉ݏ
��%
����r���M3���醭�I<T��05I\��&�S^p"V��W�~���tR��5�4
[��ϛڸi�����3k\
����l���sf95\�ͳ~�r��2(���;\�ُ�"}Vň1O�/="��oh�<E��
P��gX��e��)��[��w���*I>G	�'\3�:(a�����u���L��O菤�xە�3Ɉ��Y`�1ИqB|���H�����s2;�i vτ�Ÿ	��'�ʓ�4
ƍ��|��Bs�F�5:��,��X�$-"4��
�XRo�{�p���i��%3�;q�Mz}~bJtWi�T�,h��s�]w��0�9��w�d0#|DP�.�@F(��>��@[�� ��/GǷ���^?-\�guߑ(Pb��a�F�:�'�%Ӆj�V\�w��}��~ƾ�z�E���g�k(
��Dҹ6���7�Z�NV'�JRG\[A�MX����������"9�QހC�jf�f�jP	���TS���L�t'�/�d^��Z3�5)c�0��o`�ثQ.�m&)z+�����EWT��'{�f��;�`∮A��*{��	�F��b� �l�BJϊ���_����N��r���W��f��E�vg����&�'d�X>�.��\��"��ex�����' M�����*kpL%<H���{N!����]p�Bil�,y��1jL7r X�U�q-��g��5Uw�+�	��G�`7�d�mL��oy2��G/Z�k_���}勚Pi�mV+Ӥ�z���h��B�CE�q���q��I �����L T�����3���A�W�w9ܗ3U��������we�ӖxC,q��p�'JK��DKג#�R�d�	�$p7�C*����x���H_���z�)g�u��U�Tm����W�� �ˈ��t�/�b��$W��y�ݺ�U�r��`~ުV ��z��~��K?3�Ӣ��d�H"�Y]+�^�f�f�t������uN�.+?�Ə���{o<����@���6b:Z�ꆉ�ϭvC]��2�L����GB���E	O��u�@�סϦM$��-��4g9#ƈ����~/�즪�Q�Ū6J���q�G7W�6Ǖ�Jm2r�{�G��?�mU��Íi�8�%F�1A�V��IGQǌ-޴x�iA��+�c����FOCď{�9ۙq�D���8/��^��Nտ�m�1�����ƃ����m�
�̑r��sM�4θd�F]qy?�[k�HVz�"���k6��"q�z�d.�bD,���&�C8�M�)p;k�\�T�UTf������~Nbr�I��՝)"�<.�}Ɂ����Q0\�����6/
����R����H>ejo@���?:C<�y�#$o�!G�Csb�bs:��K�&��y+�]���8RK H.~� !Pf!����sgҎ���W�]�b����w�c{���͸���������eqϛj��x5�*d�,�68>4+
�!EҞ�ç1O�D���z�^�щ��5�BF{#v:|��؜�ˎ�w0�I���?#���� ��af�ţ��s�F	ي����%?H'���0����W�續�ru���2vpFB�|/g�ت��y��{�<�����Ȩ�x'�D����E����#HH27�N
�Tc ���G����M´	��Sv�~�d���M	*@5�u��4J63kD^����7�[j+�}w�&����
�(���k���@�&�k�U��;����/	�y�vwW3�!M|���ݍ1ŧ��{o?��:�*#-g�r��F��j�f����JR����E҃/=��¾S?8˽0�b�6g�!�oZQ��V���"jŃ�名a�-GL|pC`^�2U�f�x:`�q�`�^$����" �#�����d�q���Ģ��R��@w�~���%~YQ���D��jq2��u� j�Ac�}���=ӹi��e[Y\pTdA~|"Ɵ��1�i�LX{��pL�ԯ	Ӟz�s�+,�B7y_<���Fr�-���#��u�C�Ugj��L�Q��v���/~�-�D~i}�Y�ײ����@�U>����p��g�<7\q�o�_��g���NJ�lE�Q�4��3Y��V�{P�2R9�`x~/d/�_����q��|��y�f�!T��l�zT��ī��!�(�8�Ә;�~��{*�+��m��!e3�4~���>��uOk����Bbd	���1��z̖j���"�=5S�#����9�����8�W��.{_ ,��5��h�-��+����˛2]�}ɔ���� @44�kIO����	��Xq����J���
�f�uұh�$�d����B-K���r=��J��;���� &Wx�ďR��AC�*x񨊏�B(^ŷ�)W��hJG��B�O�ġ��]m���*d :6��qJ4�f�Q��&���;nyME���٩�b�Y �@ҭ��j�p�q�]��i�&;�M�i-��~~e�/���;YQ5�>b��CВ�qZ*7@��ݮ
� +;����pż%lC ��A{��@)�#������������Xt�C&
�(2���L�߅�D��L���o[����$Չn�1^��� ��q!��'w�J��OO�]�BL��0�f�*s��I�%cr�Q�c�m[����<Y����^�����S+���/W���x׃�O+Z~w1�@��+3�s��s'��\��ù%�gf_�ذŪ.G|D��*zEGL2�gC�ej��b�O,$�a0���FZ�ٙ9{��S�8�[���=aqr����������E����4���Z&(Uc��	��u<H�׋Ud�a/9.�}��J��p���.8������ۥ��t;��9��_b">i��S��ٟXx�36�<q�w����N��	��Ć p���/����*�^��8>cg��=��F�5��`GL2w8"d,Vr��{,8�%D��*�-K`�^�a.�('��D����U��޸=\��+g/��b�S�*����<���&��)��2�+N�TT-�
p{�{,G�O�޳Ojuc�5܇H���9WD��P�C�0I����[�Qi��Gar�oT���%�E�[p�ٓl�<b��B�7��I-�貋�|�O}�q(5"#݅?�ķ�x_�5�P��ȫt��>q���	g�m��8���!:�:�����{��MTE+���v����GQDNbpa��g"#օ��zݮ����H�A,�q�}���r`�t�pjU��QIt�N��ߤ����#3��q'qa�e���d����*o'}�~pLkpAe����3j�q)L<�_����Ķ��$��FTi���ƸBZ��k���p2��C����ȞJ�t@dM�2햰Q��"���Da�4�L�_A�I��I���^*���9en�_��C�I�J}��V�I�#���'%� ��{��bSf��)-��(R���ʐ|G����׼n�31QH�5��x�֏�c$��y��:Xfdtj;��>��39�b�q|�7;�������b�����R(�Z�D��J2��(�KD��(�܊�T���A&���bSb������a{�L�|�	a��>'�<C[JqxVb�}D©�m��ܽS��/��F}�fv��/r��L���N�Xt$/�|��ϬpQ)��`��2,��bz�GXs�$w��Є�41�.n��*�7K�o̕9ܝ?�t�I~�X=ss2��tz�P����NtӸ�S"�|Of`�.�.�M�0�N���K� �B �g����ªy�ޔ�)�7�_�+">�adÏ�9.���ղƩ���L������9g#�&6���$ ����Q�o�h�r_0���D�U�D�N.��"@�I8�J)m��u�ǭ���rqo�ܒ�jq?o�fzB��GBdՅZ@�c���h"v5��PA�$~S��^�kc��߅gX��&��:4hAp�����C��� �n��I�s���M�s��k�o�EN �����zjF�]�͹�#�4�b��ls���T�J�
�.[�g��x�pbH�B�S�X���ɽ����7C���c�k�&yw��g�o"��v{��1{͝���#YtK��mՃ/�`u���;2���ȉ\lkh9�@	ύ�ßs8X!>�j�j�$m�H%� OQm�g�7}tL����N�z
I8ɡg�i���h���	�:�Q0�0�m��Wr=�c�M>�Ey�P�#�	���j_��6O���o��\��:܁��{a���'��:�%U�°u&o�>��T-��E���M��~�$C�vk^)|���'���omJ_��|wzh��ꭔ�C^
�aH�ǋ����|C�/� q��ey��� �;�Xe�,TU�'/Dc��-�ř�8a�NIx�6��o�V����7ɧ[���[݌Vnb]�����2��X����Qsn%h��iH���02�pn�p�Ei�K�r��;̦���nG�v�@�!aA�*)�Ӑ�Ɓ�:�`��0x��f���y!b�NnĿN"�ik���F�5�3S�����OL({���C��\֫g'Q��,��H����aD`0��	�|��W�3]�,~Zu�����t�&<��J}����5MT� ^#�k�5) ��'�觤N�ޘ�y�XIA؟{q�Ur|b�W�+u��.��@j�\����ʒY8��m�W�u��1^ΐ�9�"r�W��1/S�d�� EE�$��� �J�Xkty2Z�`�S5	9U?$��k�%�LQ𦓮VD�SطQ8���Vp��*sTe-�e�����1y[
5�3y��݉�^n�xD��xZ����CV�ͫŇ��������y\�N^��
P4�4�]��V<�SH��_���xH�~��8�u���h!Z���@�!2��⣗����jeg���z�/��^�k�K�!��X�k��w�i�:�:	pvM蛚 ��*�	�?��׭��Vu�k�2�K��������PtԔ�m��޴������S��gƾ�X���f���B��t�=���>|�'{5��g6��m�G%�Ю">����!�_��J�rx\<�v�^�Mҭ	�c�w�E��A3rkeT�"W$�X�����rܪ�Xm����z�;�97ʀSEd��܅h�x���۴����� ��#h	�l+IX?�:9���;{ѫR~$��ˎW���8�F�w`�V9s���t�e~ݭ9ʩ�W\�����U�*���qR� �:��vP�t۔{8�T��@kYq
����sN�����~iu�)��������2�<E��R|�]n�9o�XN�6@��!0[/�ʙ�F �}!���ޏ��,���5�[_�U�\LV[C�Ӌ�ة�ĵ!�		kIp���ep�I
��h�������a� 3h
W�#���[����	Ju{���)^�ǿ���0����5�u:{���CC���U?Q�c�dG�rޠ6�޸�����bH8��&��3��
���7�����nbW;J'	��}�����ˇ�N)8JK��} /�>Tʻ�ձSvt�:	s� ������)o��>�X�o=��d�Բ��8�Ű�9���`�n_}�z;��*��!��;��V�	��_)�Y�d��;��&p�gޟ��vB�n����Q�9 ��	u��N��t��R��ڪߛ�f����^��Wq�Ο:� pݯ[��@@u5G�GH��v�-&b��׷Y�d5;�n#�:������{Ɵ�}�3���Q������Y}Z5��O����^N Zp�*��[Z�V��oûR���?A�fRE����s�s̞}������/��О��R	�)oH�<�ܯ:'�g t���<�G0��ı��#C�^�d��Њ�黻O�j{��;z�������"����C�gm.8՛��#◽t��{�<.j{K|΃�P�����>)���`(�e����!��tN
-��e@�ܯ�&j8c����ޮ�ؼ1��O��a�m�����\ע^qZ���p�G����jw�����  (_E�Bw���q�΄K���C��W�'���-x�y�=��{J���S
��Pؤ��>��6�V%�3�W�l����|�ޤ^���~��RB76=���D��^�����
ȃ�S�˓����e��?_F�,��Ź48�O��h�����O�"��FU�I:�I��{d��۸�=U;��@�NIw�Is]({�����ݨ��J��5C��>�|��)�����$��`Y`�AP�t��
ʇ�����@\��ot<�����u��Կ������ [�"����3�X�N��lWO�&����g6V��I���S�E.�"��O�?���G�]5��R���:!��Nub�犆\[A*ٗb�K�w���}'��l�볯�l�g�?B�����G��a�W:�o�Ђ���,�#�ጆ,u���qvꏏ�Z������h.���������q��o�����L�0\�Ɣ{���3�x��C��~���9�[_��HU	�R�ƭDx���c���Tq6��+�b����Y.GGl�sY�s� �/I-�T�-/�e�g~�އJ�O35M��f/�v�TB)>�	�+b�8xjyE&��P5;[BԜ覐Q�����Ȏ��w�v�A��A>N��8�9�T4�Wٴ��=�W��X�@Y�P#����5�J���������\#өQ���M�ʒ�t4�Վ/��P?^l���l|v� �v�J���!�$�>���q[��-�@#�戠w��6 �����<4P	Qª?w�/�G^݆Je*ۉ8y	����7��X0��=�9wj�7�=76�%t]Lrd�����-���ʗ���!Z���.�Ad�FY���C-9a(%�MK�0q���Z�ò��KN�I�c�O�K��� �io��駜+Z䵶�|17eH�o7������78�tB|>pf�e%��}�_6V��u�<F�f<�:ᨖ���������z<�P�%v�'P3w����j��f|-���r1Cտ�Y���{�����$����P�ʺ���� �>0�B6~��s�|#��Vol��鏗yu޹N˼�D÷���v��Tc����f���c�3�(*�=�F�������#�@��/�������>��~}2񌸗B��0ؕMWP��(��6�������#|���
�F���7�߸���;,�2�.�E�"˜���>\��j%7����^�4��7��.���KK������|c�
����.�F٬�`���of�O�T���=�)��0�<��K_=�e7@�J!Q�?Ƶ�����_�FI%�aG�j��:�w���v�ڧD4��E���l��&J���b���^��5j�:�w3�ǒm��_��)��"a9������8REO?����7n����V0h��l4K�X-G�m�ZYL��߹
��#'�ju|%wepp�u
�M5���r$���l�0X�����N��Z�ǂ�ጿ�����Eft�=��Hʼ��[�'��wDneq�b���yYZ��л�Г��l4X��T���wu��l#�~Z�F.��J����J:�0�$'�]
�ΗɎ�RIPU��p
m�;z�,�/W��-W��`�CK��(T�cO��Q2MJ�k�.�e^udg?��'.�qh5)I:��81Q�p����/�d���爮����C~��Z�d��?�{� Cy{��_N|h�d��N�)� a�G�)�R��Nzck��Nv8F���	S�G��z���yD5��ye�	��V���aFZ�՚�8�4�t�V�U�ڞ_)�&?,JF�EqAg�(���JX�wtT����j@x#�+ŀWc�_�,B��P$�>�,�0-����/қ��7�/s��)H��]�O�������EN�26��5�{���}	�i@�kv���o����[�2����Uơ����neMO\-Otl�OMK��/J���:T���0�ʆ��]��6�o��$�*�e����F�#�/������b���H��Y�`�lh�	��rp�W �{���]2��~ˠ{r<ҿ�h����k��wp�����}Q��1�4����Fdp��Gl�{9w�j�`D�j��9>�}20[#��L��9��w�N>9懷�?�p��'Z���������f���S�GW3��"
�>Jf�M^��y��n�9b٧\�ֺ�݂�aϦx|6}
g���#9�b	�S5��`� r݀'�\��eb]!��v�0���uc�S������s�AM>��,�bK�|�=����n�k��u��[�0��P}8a�7!��a�~��o��9c��6��Y�}�f+Pb����������O������O6wS��i-3K�\�_V�~}J�j9��gj�sS�xxM��9���g_
kO	,�]6:B���T�iس��E��*���'�'��0�Q�
Ia���g��ƞ�� :��
tߠ{:�p�4Ĩ�Ά�(�	ޛ)&Ѻq�[S��Kسl�\a�7a���ݠzT���V���q(��E+_���=�`U����H�GW�Ѩ� �ҝ��L����6�`y�/���!��r	
TEǹ;5F�4��͊�ln���ܼ��E0/�݋������{ֶ:�D�~��D�q<-�=���:�%��8�<�U�o��Q;�X��g�t����l�Q�+h��y2(٥c�}���	�F������7�ڃ���$�o5��2^��%M3�9p���@<��D�uA���.7�K'8�( !|6k��BS��\8^�'{��p��Q蓸�n������R)v���1�˩��߅}	~�6�7n%5.1�L�Ǐ��;%
ц�ʞ0--��k�Z������ �/"�M�Ȩ`	�T���27\7�>��%w8׀���]�&���[lR�keߚ��'�����2�M���hd��P�(�ٜ�uO��j�AG9G`��u�B�kO-���F䅤�B�\��Lyճ%�O�E_Vf�}j�Qpj�_��/c���߈�&�Te&!�=��*��M�`�v�<U�ƽp�tth��u��T2��3]aL������=�R�?�K�5`{Y6���C���aA��чF��qHq�)�U��L�9>^~��5�
Pou�-��_��t]�e�)p�t�*]�Kq�z�ѧL?]�C�"�T��=-���CIR��N�]������)�u�7�t����p�lI��1�y�,ͺ�Zs]&�N�I���)eUC�S{{�bˈd��e/Z�AD��W��J��3�I�H�j��/����"ӝ�wK
�:���6r��H���l��u��Lk2���#�jEN�C?U��ᙒg��u���F�.
�O�,nBt}��9z	�)��l9�sўZ���<
��*�q9 �9l���/z��h��n�A���t��������6$y��A�J�Q3��P��bT��u-��'��q�Ki����J/�m����V\�~��a���c$}JS�r�J�觴�N(US��CQ���:m#�����MC�]��bQ�n��"ʟ4v���O;rLH�x�u������R`�e�`K��֗�.{��z\<el?_q�x��s�R�P�T�zZ��ޟ���~��)�'��z�!A �$����֭��ޠ�h�R�|���չ�&$5���UhE"��5e�b/CJ���=�'�9�G��������%�����Le~���W�ښ'�H�4����v��]:���E%����kz�,���ZR����o�ֿj<( q�p��G���uò�R(�8�I��i�]#Y�aDR"�IyG�.��|�6��X���8/�O��\lB��U[c0?U*ʈ;��
u����'�]ؚ#T��կF�Ķ(�uٳ[\��Ɖ��A��!.�i(�#<�e�������}�OʱPDJ�Cb�y�S$�0���B@*�`E��N��B�Mj֌�}����?~��W�LK���:��y����pm�Ҍ��9)����5H1bo��С��<Il�X�5�����
�����L&]B�r�7R��z�	�O�h�pk?�4���IN�nAN�ꍅf>
���*#<x�@��������u��㦎�1r|�̟J�>�bp+$�`��Ge,د��7���>�"�?�f�+�T�F^.�2S�w�:�/�Qi��e��M�W���g8�y}ɜO�X��1��4Exrz2r�(����(�	�:̮��������+غ���QkLy�D��VKXLN��RGs���QV���b�@�I�:�O��CPo�ƯE��gP�z��F����_����\+m�@c{��̚�9;�I[�u�^7��N�X&� �,���N��������zX��@�a������`N��`��9��b�G�-q�E%�+��f�wG[�'X��n���
jf\x~2Dc/W����5[�~�W��e�7��0i Abc�p!�ɮBT��`�t�i��W�ɭbw�;�:�Qjt�j�z=� ����lV�6C����AN]��dU*���V�TI�S�0�k �r����JU�2��-gjQ��'��M��E�W�<J��n�wNN��Q��w�4��H3%e����r���ۨ������iP�p�0����Dղ���g�C��ê/�F�( �ffA`�A��k�#5�
u��\�s#O�3 �T5)�˱	?�^K �2Yb�`s�0u��]��T�\�cV��D#��(�-����>:���J]t## �杪"�� �&Hv�Q`���L����&�}(F�2$�g���F:��Q�6�D�JGRb�w�w�Yɝ��1�9�W�ݚ�$��L��f�Jw~}��qY�{�QWQ#��)r�,��꤬�~>���
ҁO�n���Z��,�Cީ���U�|�����J�]EG�X2n�����Ž�1��Fܑ��o�i���4��"س�g�q�P�X&_(%rrO�1������C�k�ɖ�<�V�?�iB��^�-� �8�n��":7Y���>��`�عa