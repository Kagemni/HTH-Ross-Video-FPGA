��/  �k��~1�8���~A&ɀPb�	*�z%�a:mTt���NJ.�~��uW#�i:ҽ�����=��ď�^]K|��"I'��=A�.�\߰��Yx�����7� �c�i��xWx�{�gF�6[�n����&�[����a��ʈ�
��w� ��W|֥�nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n�W��ߌN��5=�8�:N|���gp�P�ظ��U��)�& g�J����[��kxO{F�ض�����F��T���n#'ڄ��e���7��ѻ�t����+�<�g+C��H��X̱fT��%5��*����U��V�է�b��?��ڪ���Od_
�g֏�[�%mq��>�[�!z��^�,
*v��%�n<+D�';01�b��W���fx�w��SE`Q*�_�}J�I�Ff�C]�&7G�Kp�S�I=�ĎLi�.W��z��8��\���ǋ���vQ��hv�D]��i��N�@���g:d�mUGoj��'e����U7k4r��Kg�9h@��cd��I]����6�q(�s��Ae�Gs��ro��x�2��S�S�.�����N`,_W�����7�R�!m���g��}]����M�n! -qȋ�M;
g��`�V[�&C�������8 K� �J�n��̑���������<�+TQ��/�q~F���`70���ҳ�ԡ×˞Rp�h�q�Ph&��.���Y��z�- ��`�̫V�_c3K�z�}WR��x{n�W�C��X�����{NK��^.�A����cڦ$��a���+��G2��Z3�.�LUG7>�p��(B+h|���ٳ�%U�a� W;`c����\y?�io��ᎇ�f���|�_-%_�
��� h�l1�H:�ɏ��A�釀�p<*��#i�7s[k�y_	'��Ȫ��ـ����Ә��	�i�������hͳ�qʱ�p�|n�P�o��;��i1k/�����r�wt�w����,��[���7���	4	j�RY I�M
K�sH�G~*v��&��+�
�x{s�0��ֈ���%;D���N����Q�b�)��Qn�ԯۢ�Q�����T���������&k��[�	D��#;dc��8ZU}
�����[Bk�����5�K�nh��/򄚖��f����ӝ�&d!Ãu��\�v�B�<3�O�,g���gw��9.��*��G��P\�k)���ܧts5�D#1�s���Z��$��(�S.��y&��"�P��,�l�B��e?�K���*�S���F�H|�P2�^5̏��%a���37Ѡ_'�Q+�sŰ�k��)��41ύc����F�|V�T]wC@��7h<�ʤ�]��T�ztA�-�@_PZN�K�P١܌�m|����jj��
t�L凔]@��C��n4K�N� _�)t7s�>#�iG�{.�-wNl��,|�ƳQ-2-LNT�bvq�g>O�>�1�p�������$���1/��a{Kb
џM}#E���+̖c����&���ފ�nH=���,v���;��6n���Q�:���	l	_i��,\2K���K�����)>=�r�8����e�Sd̜i��%��:�/�I�:Α��G���<�l���<F	��VjP���|�{�=����$�+A��{��:�l�����'��Ẹ�x [���Q.��9 M}��˷#z~��v��;���!�>�aּWuG���!������8ΐE�͏8̪�|&7@����+f�@V8�����Y�m��\p��2�t(Hpk5q�����/ON���������
ǹ'�2���/�Jy"�~E�5���<���D@a�N	�XFO��R���Gf�����I��0��<.����7fKo"ę��pɧk�nVidG��@���^����w��P"�16Iv�P�?��y�|i9�O�k����r���Q�3/�� -�-X�"��Q9n3Aa<W�t0)H�
r/-��Q�4��Z���b�bUz�̧�~noѻtM��߬�ؘ�,319�S����/n֖]����v�?���-t��i�9S�}~���e�9Ykv��O\H�|����G8�����f���5:]M��.�.0�0_tG���ގ��~�$��<�8g5Ğ
��_���e�R�
`h�H���Z�x�z�F�r����D��cc��]�\��'~�I�z�`�b��2��[j[����۠if�?{�bz̹�h�	��rn�D�T�:�Zt���AJ���ӯU��>�0��O���0�h�9)�j�o6�,��o�z@;G���!���9T	
 ]#� ���y�w�<u _�[�9*�s(�Za�)zF�6�~��3
m5�vd~	�����|���t�w��� �=Wu^w(`x�@�\�t�!?��{j���[ܺ���/-@�� ݙ�H&ȣ�ɻi���ǉv�}-=�?�bOr?L�B~RBQI��X�"q#���v��3����di���R�ڤ�p;���Q����\��g���*�'X�B3�h�k�;@K�����7o0�	������~X���󛷜������*���=��_�=ju-^�A�`�-�))��d)�P�&fV�~��"u��<�	>�|�� ?��Q��U�ڕ�4����V3��6К��`��̈[PEf�+��l&,]8������ت��������ͩ���)B�,��3��G.��t�v��0`�*�I Rj������ �b�6��������Q�B_�[�>$6��{O�ݭ����/��o�r6�pgl^�w��^���������-0���e����_,��t_&�:T��<fC�oP��7؂��Ô~����!|�?�i��t�|�PS���NU���IJ�;]U<��6*�>u���_+1� մ�n�XbV��n�ˢ�'W�n�{{��\����cB)d"�}�B�q�ʹ�b��P1�!��cB��Gbq��Ļs�o1�1'37Ҫѷ�vi�&D��2���V8d�"d��L�A3ށ����b�b�;�.�c"��i�r!'E=������Le
�F7X�Oy�0Y�e3ꎎ�GYn�xeX4��-
���
.3DX���pD�[��o{޽�
wZ�w~!���;�1r��Bs�;N`�����C���^Z�m1SP�v��ej��i�J��;��>~#Hup¹�ByJ=�)�!�%�r5���|�^���1�<_8YAހ#fH+��D� ���d��ʿB�xb�5h���>s��K��BM^����$%�q^�Ӯ�FG�`ϯ(��7v4��vśi[��^S�7i�J�M��5��65h�c2n��TѺ����5+"�B�Ѽ�'i޾��<��4�M��9��;Ą !GheLm�������BI�4�q\
��սxm�IJS�|�|��줐���$�G%`Ҥ+�$���<h�v1(�ZT�s*���KX�_ڬ-�Z�����0�RA'�>�6-��)fmhî���
��ߧ*6��_�A���@C� �� �*;�0+��5[��`k�[X�z-]�.5����?H�����@��7��1����t�D �ouBJ+�.��*Tgk�b�-Sk��zE�0���2�Eqk�FE6�Ӱ�,eN9?x��`��) ��QN��n!WbU`����m"�ŏ�/������6s`)����F0R�Mpv���wT�K6N�&S?���{� �z�5�Bpͪ_�N_�Կ1�Ƽ^2\�����<�����b��^�P��vB���$^|S��UѦD�kţ.N���ٍ�Y�)}0B��6�_�NZ�.d~��`��]���W��]�i�I��1����{�>����%G�%�(b2FBCݯ�g
��x�BR���:ö &.��Ҝ���� ʃ6�T�E����^��	hsR���^���,p��M$n$�ِ��bn��/)�첟��H�
���I� ��Z:���r�ϽM"��5FB��]������0[�#�H�r�H�~�Wa��Y�w޽��-������p 3[(�Q畕[����
����+N7�pe�4V�_��k
�ŉ@�,ܜ���f�9�|=��٭L�`8���(� �W��ռBm����a� �w�.��z[	�ě������d�����W"���>��JwW�i�R<���ƥ^ �Nd�r��#��g�wÐ]����I��ER=�$(��Z%*�`D2�8L-��	����;���%/�r��UcM�JMRi*�T>��#b�W���P��X�����Fʓ���\��;�w'Z_�&�l�����n��k\���b��cY��� ����}�dո�-&x
�"�H!/E[�<��T%'"ێWWL��U�L�(A�J�K���U�� �4����U�e��6��T''���^�Y��mh��cL g�Y���Ʋ% ���ٌr�� �?CPGL�}w��$��� ]��ʿ�?n9Ԙ�R(LD,ϣO�Oe�� ���"����D}��� GV��|����:��b=�R�rH?9kf���~��9=�����m���1u$�	(�0��&�h�
���8E�x�*%����3�RU^Uz���a�dB��h��T�w�D&4�3h�}\DY��x�;��[�7|�9M�Q�M;��n��-U�9��y��{EP��@M�ɹ{���[�('�j�7W��=�C�ko�ܡ��ֺ��!�S���WP<$�i��#`w67^�!�
��4��o^1�S�I�q��^����Ct�
7p�늕v"t�l4�T1p�°pj��j(,��X3��_�t��{�x ��٥@?~Xp6E��Df&\���d���8�"Qj,��$]�3�=i$%�t�ө$��3Q�$�D�WQ�Ė�`y&�g��(^4���r{5��I�Yڙ���Ƭ4(;�8���J�(^�S�B�fgRij&^�V�x�l�������~DV�ֵP�m�gt� KEÆ�������}�M�F�ԉ�W��S%;[>�r��Sh����;=>���\s�	8��u1��ޑ������[��e)u��"���)"�O��l���V����u���pB�Y��=~��u|�ח�hDZ��us�w��UW 9r�	P����i|�P��Gȫ������L��h��n������3�>gd����3*,� mws�R��{��������IL``P�^0'��c~@S7G(������wn+m^(@�Man���0���۾���F@/[XcJ�I���ɐ$�!D?���;2d$7���@@*J�*�霿p��g�)�6K�'�hC��IZ�.	�C��%(DM��h���)z��Ӿ=X���`S�ܼ����P�S�L��ℐzJri�B�(��ԲX�����$�'u���]v�r�,�\�6����~����E�:~�r,hɈ&��Q�>^\�������4��ž����L1cׄ����W�8V"�HF�С���0��1X<f-��aXK&�~�*^�9S{��3�ֿs$�4#
�"4 �� �\�JBNv��l�IHT��W�*��|D�ʸ�:b�rʦ�*��e(�C�r*����<⅀/����B|��>$+�v�8#�ވ��uӵ�O��w�N�ԣk ��3g?<7jD�?ϛ��+����r�ZE�V����)�ꚙg�k�=��j��j\� ��ܰGx!>m�#FJ��y8�n�X���E��y6ǚh|(l?V��e���pRM��7�ɸf�.�"ǥ����+�V� �MB��������%!���:A!��l��mc�\��>�s�r�̱���N�Q�vҤ6!�(쒴��cU����3�~{^ն��N�R���vC�6�K5ڡl��S������D�W������q�ԕ�~�S��웛̄
W�ф���6�Vs�;G-�����(��X���O��R��S�No����2=q�O8xn4q&'�p�)�fW���T���J���_�s�c�MF��%����=\8_������.4[Wf�2����W���/��\�E���Mqn��5I�n��my�*b-oB��t*зe��$��ٿ����{C���j�H�3�Ur� �QC��PEj�F�D5�&�>�kB�e�����,S���=�]��*�Ik�V2h-�!�RX�Jsf�{hct�2L�A�ǝ ���%1�7�EK |t�[ ʴ�ss�j��fƍC)~������~2i�t޾]��(�8���@�	�	���6��������q�N��rm�50�0�]pD�@�Ⱥ�����W4E=��:�!�*g������7E"fR}Ņ>�ԛ�ȑ� �m��.y{	���"�	��QsdI�=�m�
̦�o�+q8LR��a����\��ƨܮ���Y����@\���q�e]�А��ar�	�u= 07X�7�|/="5
���G�!b�?͠���a���7~�l�h�gc�h�*�ԐFUS/�pc5A4&��6z�"|����_��~s"~����k���?)JDZ��-N[���ٍ�Н�-���������^ ���"���#������JpDy�#l�3ע1`�:�h�0���\V�V�W"b�1�Z��- ��T��^�ҹ�(�Mvn��,(Z%�~j_��jY��w�Z]��3N�Rz��E�-��w�F/t�����������@ay�V�'�	LTV�|w��j����bc4f��]kV����&�,�է�oܭ���2^^ȿ���L-��9�_b�+�]�Tu�ӓ![r��Ɠg����~@�Tש�ɰ��(u.��s	R����y�v�v!>��8u��.�dŔ��1 �u4Q�R��	�8��ǍIѨ?^��'�} ��0�\�7�)�����Bh2��2@~�HD��}�7�����n�R��h�>G�a��Q �!_�aD��Ft���6+mG�Ԋ��m�d����� �_K��U�$�N��|>d�9�%X8�o����'���I��>���jF�@;�]Q�J�ғ�o���[�3qT�J|�����&��@�J��|~�b�����C���㴴�)0SX��	����j�Ѕ8+��W�2lM�_�X#�Y�0�F������7�8��`%��,-�6�_ϋ�h^Q����c�#P������s�W�V"�j�����6�Cj8<\��@͇)|b���>�A�3Խ�Z����-��6Hق�р3\TJ���(	��r���8q��S`&����V3S!�-�\���oҶ7$��1ل�.���ͼ\���h�����,G��0��s ��Q
�ȴ��W��h~�v���߈ԑ,�������E��<�>}���^���,�?�-W8��cCP�cH��B�)�A�̲����z�N��V�����V���sZt�_� n�q�����WU��T����t &����{�c��QV��z���-α��%��;��w'��
h�\�0jw#��O�ce��_Mo�)G)���}��Ҋa���T�{�%��*<8����#r��F�r��Prp�pPUQV�l�>G�w-��պ@�Ku�^���;�w.�&�f!��V�i�d�_яYr��x��sfb���#��T*���b�T���<GAxc�>�[��.���~m��i��I:e�m�	���y����pȓ*�v��ҟ�4]��x�G��ck2�۞���~d�$S�k߈o�@�%9	��Ifx	O�O����#���&�������F�JG}8Ȑ�����C�0n��P@�o��l���Dlڸ�^o3ն��xs8��8:2��960�l)����`cP�1�~��<�t6��.�
O�zV�mC�b��<�7�FS�˸}/�'^}U ʺ��܆�rS���1���[I��x�߂�c��rYG�F�p�s�����a�x���X�r�g��Ә��'�+!����O��W�"X��#��M��d�����
���Mq��q�2)\,��x`��wͬ��ǀR;��!�[���
�(�/�J?�0?�v1F�H(��A�)�nz̸f���pA1}u��W�lr<4��~�f�3�pg�챕��1gԬ2�Z�*6ITm��7$�88M;�Jc����-����I�H4��%���(9�.�t=�����ޑ)�����(����h{��=��UR�������cn��@�}d�(��:u<�A��r�����(gP������t-qf�����Ԍu�oY�O�3D���T�keC�����4�DG�Ǽf�IS ����Ϣa����[�_��(B�e��U��޲Ɉ�G� �N�h�h �c��k]�ȷQ�RH�\	�^��	�x>���:�)ˏN�T�r*�B�[/�9�\e�aHYg����0�T�B a"���T!�(ʰp�/=&�� 