��/  ��0^����I�X{՘:�,RYM�r�4�����|�|l%��4�<Φ���Oy���I���g[�O�"`��S9�I�%Ŝ�P���'�����t���T���H�n��+�WN��j��*"w���T���X�ǳ%h�&��iqu�$e��s ۥ�nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n�||�p1��b<o0]�z��L�^6'
I�B��������"z�S���')y��oK�W�xZj� ��r�m�χ��ݝ�S��ݤv՜+�⧩̙;4�ܼ)�9�~#�@�7�K\z�ӊ�%Ey��Ũ��i��{���eAZ=���ަ���N���.�7��l��1,G`v"�z7��J�3&�yLՉs�2_���K*R��@�^��e4��僇����������B4�T������B���_��.�Lxԯ@<?�p�[�|�T���mB}���Ĵɷ����ժ+*.��}�a�z&*O��h���u�~߭yJ����V��zQ������;R�ӃkyX	�E���ܚ�Wt��H�;�����E"���3
cw�]�~�t�i��[6+��h�n2�H�:����x��B�Ԁ�+y^a�R�+�O搲:-#k��l�w��}�����t3y�L�:y�C>�]hT]�R�����T5�`�$��d>뇜n<�/����T��N��%��c$�͗zN�T��s$n^?��*e�������dnx�hƍ!`�8�
-{�'��1�C�ᨳS���/�/
�a�آo�Ե�^}�����I�cnt�G�|Y��`�^�Lle�s}	�tP�u:�9J�l5��>���6V'٢��^����#�ɯ|3I�ڤ�.�>\�{Q������f��v�����-�E8P=���;+D��7dA��F�tNzf�?9-����P���������u�m뙢�29�x�z1�|��d�I�׫ESܫ�a��D�]��d�90���~WMh?E��S_�FL2⋆:D-Ja�4��0J~�߹��+f]����ou�D����Ѝ��g$���ր9@�7v�hO��8� ������.f��g�շ�I��ĉ|������B����(N?��'EP����b�c�0�')�  }�m$J�R����0Sf^�T'�%	�,�,��-�0M�$� ���+ONp~Ɖ|�����#P�~�ښ4�+�D�����Z��v�!�5؅�J/}7H/�*I9���?������NUH�F+� Ifk�`i�9[�;��ʜ7�L1�nd������pK�F��Jn�T��`	��ȸ-�Tj�Ҽ;�9�Z�^\�b=����e|�.嫸H��zj%a\�|�T�?˥)Фx�Z��*M�6>
��s�Ơ;������<C�p��s%�$U�+�^��;��U���k_�&Y�D�g����*F�i���0e��J���vbT⫞�|�����1�3�ʦ��e9��m�����@k��v�����(/���|F�.!��+T'�`�x-gg���}I�:�v�	}�iG�k�lڷ�5����<���c�;؇��F����V��͙'-[4q��	���|L�@�A�ymvs���N�\��H��1�1,�p/���ވ�*�5{��=��a�z$��d�@���TK�C^d���o�S<���e�	��zЗ΍�T�X�vW���a{�,\!L��t�p���&y8�Q�/^�O�r��@�Il臋��ٱ`��+�vMq�B�~�q#2����D^�V����1�L���⻗pIWQqlr&^���3��^ �S{
�,-�æ|�s��!�t�J��%�8�U��r����|�RB�y�~"�|���e��ϧ�n_�_�2_�g<2-��y(��]�ŷ.�R1E�xj�㚲����R�{F�.D	�ۂ����NW�g˳1*�(.��"fB���W&�6lFfE��%1|$�m�泑*��P���g������'�Cǃ����0'C<n�LR�F�yvS�T{�5����Mz��y��uҪ�͘��E���3��V餯_:��nKt㔳EF5Q-�إr��J�5G��!�By��D{��Cj�.����]C�ǜ{gy����No��9�S"�P�Mwī�����,�~����MOX@�H��}θ6��-�ocB��>��!�W��:i�2�!��������:�D�R�<B���xW�m�tߒ�ZTWט����;���`�v>���|8]ݥNķ��� ���ߞT�@���/X@wu-�Mz���b��cx�P&i�o4$�Q*�P^�_���O��tI��iv�,���(x���}SU���`jO���5=���x��̦[zw����K����ΝG)��
�gI� ]x��6�E'"<����n�����ӛ��7voX7�/(��e�g��z��;����>r���.U������%)��B������G"9<�8����~.���p�i��<������V��r�R��I�:Y�M�_:O��)����.�4����B$�d�� �����j�z�a�!����"����ɔ�;+A�s3�=�:H��ozI�ԯ��]r�ub_�eL��:�J���7�d�&���W,��/*���7�ʭ�W;��Iv���ml�h�_�����"��̜6a�}�n��Qi^�?��MhE��m�R��;�U@	`Q��iL�. ��R9�X)P��O�/��)����5;�i�&�=�~TŃ�^e�HT���+���ߓx� ]ՠO	J;עĢZ����@�@�f���F�(�r�@�w�R���V} �����m1�ɬ{Z7TN=�78������0�����c��j�%ϼ�} �"�F���
�u� �9�G��y��!D��Q1b*��#ޢՅoC��C��j�ZN h��d<���)����3=���H�mV��m�f�����IqcՋ2�su�Ruo +g�WB9��������n�mj�f��UN���(v�D�ۚL,�n�Θ����f���7���يG
�-��Λ�_Y2�iݎ�T�]�X��-�[r�B���!�}�����S쏜{���B��X����q�BB"�;�.�Q��M���6��F�P�'�~�� F}�H�o��m������Qi�NaB�E�u���Z/yD�QY��3�ZZȚ�<%Ad��%�:8&��̼Ǘ�$Ţ��z�I=���SNuTE�,+b"��oc��חZ�H&�L����F�^�KPB��Y�"u���,��ݪRl]~|G�].|(���ܕ�x?Ρ�5$�b|��uL�kbMEf��xL���!xO =@vN��C��F�/�֕����lk�Eb�B��:�bʿ(���|���N�+a�����c�����W٣꺚��zBG���x��f����eSO�(�l�v�lM�F�E�آ WZ�@Y@3�����z�а�����%�/�9,#/vT�I��O8B^f����jW�:X)�% е�����lz�Lƥ�<����g�^��Ǫ��%Լ�|��(��x5��˪L�o�`8��!��mYg��OEe]5'���.��l8���6�m{�_��Y����#|t(\�)��Ի%�V�p��cO�}�dP6���%>S����z�|�.��mKx��W%�Z��e��-G�~K�=��ҁi?�4f���%�ア�����|c�^����Ko,�C,3�d]��	V�>�L�;�b�"Z��fiǋ����JP��	�˰���i��0U1�1�pٙ�4�.8�Ӳ1�Bb��o϶�Q3��*��*�8��C
�nοFۨ�e