��/  /ő؎��>�"c��K}#�h}D,��� W���G���B�;$��ʀi��B��A������c�S��@�^xC��.���r������Y?������σ9�C����bX�U���c]�ݮal|�����՟��7�9ӍKaǫ��$��]�ѥ�nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n�W��ߌN��5=�8�:N|���gp�P�ظ��U��)�& g�J����[��kC���Rm�=�����)V*�;���q�`��:vCp+���$�m֌�2N�+�s�H��};ֈo�������$MRm���1�op��5XX��
@x�o=�dZ���mH�x�N��P�_�n)��SC�NZcU���fj����@�Ш�-KV��Ot�*�����������(�D"X�_���70����X��? �䰰9d���d%YV
�fi���Z� �#7+��*�(�إF�d����Av���왌%���	��#�~E;v���>�咸�^u�
��zM̫>�[8��Oce�>N:p�t��θ���fG���17R5Z�l�� ?���ߤ��q�?Gvd�5kM�2@	+h����d<>+*�O����;���q8�V�1۸5��p'�0bӚ�7��g���A���Rzl�$xwE�{,�V�%�P����V9�u�7�t4�9^+�N��JVD�*e7���F����������C��(1��=�� E6�0��AKP���˒��{8XL�k�F^����G�����t�����˷i=�T�̥�����*��B�PmR\�X^*�Dr�=�>�Y�?�)�BE5��Xf�H�ghz+�<��?ȿ������O,k��7#D�'iܺ��pN��A��>�9�uN�FUG��%P �ʰ��k�|fI:�����_��Ф�i�g༙�I;u]L���د��N;I��__��,'����Q����e�c
�' ˠ���ٺ��鱄�{�j��_|�T*	�<����+���
{ �`�Ձ�a��"�z���Q�E�L�A�:~����$˘��-[�f��dR>��3�g�Ȥk�5O�_���C��J�EQ1���Q.,�
�1#]fO��ӭ����DY�Z�rܞ����>"���t"�4O>0k��̧��M�K؊���i���&�Y��D�ia�Y����c!�7��n	�H5s"�,��Ul�|�)~��s��~U#z0O-u�91Kޑy��l����8��$}|��!4�%��1.�Gʍ�� �l�����;_��2o��>7��[z�^��}M�|�Vj���"Ut�SLW��2	�;�&{�xK��߉D�S7dr��1��7���&7c��c��%�S���;]�"�Qv� f��n��d*vɛ�cS�R璶��:�N����%�ច�Z��؋%4�V{7��x�	*�y��*�q��ڗ^�Ri}b��I,��+ܯH�[�e�Q�`�����r�_���8(ި| 2��T^��Q��d*^ɺ�A�  $��i#��Tz�d�F�_�+R̵|�G�u�Ē���k�����f�E_��jR�{s�mԄ��:�P��m���y4�a��:�K��Yc���e�_7��h��RW_����$�5;�6&��lDe��j ��ҳO��ap5����˿[����y�
?�)S��V�ܶ�Bh��][_�,<v����Q�
ՠ�Dz#�Y�oVt�l��j$M
�"��+%ƣ��* -}�B�Ĺ�5*��Gz�G���!V�6�"���u��y{�*��ٷXr���8�B�6E�Z�;YTm��.�$���4���eU'u��=��1T!ǀ�=�-�������C#M���̚�o^��,S��&#�@$���2��,��WO�)������0�ha���vu�bb�Yb��u{���D����G����7����*|	��e���6�� ����h���u�ث�_k��Xη����2!��V9y!h��W!D�F���v�{�G�h�KJe��cݥ@�E�;rO(=LR`œ˚q.�s!��yW2L6�*Y	���{᳡��_~+{<�}l��,���Pe�Gs��9��Z���F���>'h���Έ>פm�oп��)W|\���bAk	���Ǌ>�P#�X�̵ h�0s����Ĭej���f��H����ƪ�t:���e�B��xh��bfK���-(�ծg,E�����/�� �(�Ӫ�Y:�s�n�,Xc�	�k�.>l��md\�7���I�koY��޽0�Mq�I��~�GU1+�"�0�����哗9u�O����P�t���
��z�/j�b��Um<e�g����Iq�j��P��B�,��&�'3)�4��J���l;�qJ_���]�O_��_�I�,�Y% O.:�~/���S�����H�U���7������É��"��nT��{Dt�+����7"�Ⱃ�	/�
o��ݑ����Qo~�CD)�e���*T��sE2D��*�W��%��"�X(�`Ԯ��>���և��hŷG&�W��'T<8i;�b�5�DCl��Y�^��g��j��J`1�`/�hQ��T/'���L�0��Hܟ�_�Rz`��G5�-z',p:W��9�p�ǓBZ�m���'/{~��0�Q#��^y���ר�}���8���L�#�Țm|5��!�?/��?��-�1�E3�]�x�;M'&d/�sq�uXL]�6�������v�
���78��"K|@ڧ>NH����/�LW&~
�߲\Q,���!լ���w��{�x�mD���:۪�j�U}�6_��Z�P�����Á	7Kϟ���� g
�i�	�dZ�QJD�����9}:��D�kV*ui�w�,�w��DuZ�g�2W�^:�x<�C����=M%��x�M����*�b��$��t���E\�TiJm������σBao���G�ç��g�(@��@�m��>��j#�d<�vn�>/�5ߧ�i��t'�;/�7���^NC��qJ�U�C�F�vL��4��9G�s�D�X\�h���ɪT�DMҖ�u��f�L�N�4<�`Y*�!h���GI<h&L���S��e�P�$C��<(�l�p le:�fA�x��Aلuy�`�L���EY.�f��th�#R� !�[mg�R���0oF�n醽�.��TR9bM';�j�f?/�l�"�H�s3*G�	�zO솅��%\=B������; �)Rs=��Y2bW�V$�D(���7S}�s��*�E]z
Օs�K�O��UX�y3}Ml�̙������k:ó��:�R	���h#e��i;�pk�|��%�	�w�Dq'��@52�?��wĭγyy&��J@q�T�7�=���
��}��]V�F����@ۄ�m����$��4��]�2
	7n1E�D�5F����~X��2�^t�,dWƵ 8�+�_Nb��Ko���5���&�i�5��,�%	5S����-8��c����wȷ�,��E�34"�m��4S)=y���·�Ukטu�Y��Ed,$K��� ��%F���� 	E��m��ª�p�`��ǥj\Ż���o���}|��b��@ *�MN/r���,,���'�����Iǁ(�����0~�eIZ?��:]i�R�`T��4��<�l=h~�Pj�!�C�뭬���J�zb���zF�*܏G�Uʊ�S�aW7F�@�|�&	�ٵB��[��V�2����J��.�[@�52x*n�V���}�w#�����F�Yؤ�_+R4��r�#�q��]y_�H!��V=,�{/�kfa�#�.eHY^Q�2�T[�q���;���T>������W�����s���#L7<x�2�|T��S�0Tϗ�jNޚ������w�܉~1���&�����a\����)f[�������r�������1�	�(��wڅ4��3|R��9��yA`B�F�m��·g4+����A�yDz��rA7�E1�~�.]�#/ӣl�.�#p��-���:����f��.)H�zϟ��;ϧ����+Ӹ.�[^�/#F9�>�k[�d��4���Mi'�/�i=~�O�6	~���y�Á���2��4Jj���ȣ=u�Ȗ��Wh�an�=���}��?Ly��b���z��V[ډ�>��g�T��S����ڸ�A\�O����j�̛��z��M��jG�¸�j���SС���n}k�ERB`��nx6�?�q�ۢd%;��V�5�e��+,Zӌ��1Z���ߗ�a&
	%��WCbqn��dK#��N6&b�.�T1�\��V��Y��:�$i�
��E�&�n���TP2��,�?�6�����o�J��d9��4��w��ᒕ�$�������[;t���O�6Nv:����3K;u8�9D"�'}N����q����Dw���fF����۽�VC����<J��;Ҫ���^5#�"��Pŉ������yt��A+f�;�"z��}�?��;���2kV��]�,�o��ԡW�C\�=`B^�ǫo�!�����ESS�l�޻bh�{�@Su �M���D������֤��%;��U�r,w�C��{Y|f�ujU�.���fg���9|��jf��TjGg����x�v��P5�Jщ\����h�/(�C]��Y&�X��/�~;z��>��:Q��zjP�����H��pG���C��'��*q�g�3��㭁����/N�ٴ��C�o�5�le3����tA�?�\��o�3fgq�#�Kf_Qh�t���R«��p��'�ΐ�+�p�zz���E���iõS���\�1](n�A(��� _���#��Z;�)��<�DdW_l0�`��e�� X�C]�n�����X�(E�p	"�ǃQ�F��Uf��H���yv[�~�|Q		 	\�7���4��x�p��#$��ՙ�1�S*�E�u;���<!�� ͆e�_�v�b�A�uW�)D��N{!��T���P:r�Sϸ8��v��q�[�gu��EFk�pN�׋�{�?�M��$��x�[�)3��a^hڶ =}̜X�t���m��ϣ����!�.�)��<H�s��l9>.B8dl��*��~��U�Zj��Mr�<c`(F�}�b �s�1^k	�a��x�n��1����5�0R��¬�H'�ʠO!>�S
^|$P ��L�L<��sF0�:)U�g��SC�����SE��P-���A%�J8�.��HgV_����ؕNQ�U�kQgCy��&�,�.JH�j����m �6��~�';9x��/�H2�U�G��)n��#w;������ 4��s0������=�љ�q7@����O`��X�۔�Vn�QBܐR��wn���7VB>����Z\���� qgU��>���}����LK�WH�a-A�ҥhx�+Iy�r���cfMܟ�D�u���wO$�{�.q��i��[���+�>*�Yg���t��(Ptq�7�9�A��]M�q�^R#����}E\ _��dQ�.�VB���=�D���>��ʶ��ʓH�C��ꂗ\�xm}��L�)�h��M'�!�m�$^���1��*��#�bj>�T�Jx{��#@֑q�H�,q`�b�[�?�-��K��A��)��4����w*���Xb�e>��ϥ8��߷`vF������\,r�� �}��Q��0���A���/���=�kg���ڕrCj޵���W2���Z��ΟR��-�y�Ib^�	Ե=�'fHùs� �9&�eϏ�p����������`KH������� '
��4@UvYE�����z0l*���PPXO�gIա���F��j-��#��^�g�0˻_���b{	>���ʃi�����3��w�j�)���R���ݛr��Js�������D����_�a<j��ż ?�'-���	�ז^�ɝ���@��l�K�;l1� ���.��KĞ�u�x3q��f٣#(o�Ǜ��I�ڤ��A7��|��efs�Ê� "6�(��Vt�w5��u �nOi�4�.�Zn�W��V�wF�����(||�{b*�Ȏh�����i�~��`�;xa� ��������E�z��4;2�uSr~�I� z�S�[�:j� �`R�x�*:�ra"�v)�\�=L�1�=m�Y� [�y@��a�"�'х?X�	Դº�:�k�� ��f�WO�|)�D���}��GK�bF����2ZpPw���F������F�M	~�V}�H1��0��x�q*�u!hp	�,0�%��</Z�6X?��Ձ� �[�F��u���*Q�6����X�ި�����~>Ώ2� �)*i�Y*R�����|u�������ݻK��x6Om����ټF��F|�EP?���=��@��.x
���H��Ï��{w�{�ߢ��r@x;*�z3����K���Oo7���>��y@ͷ��w8t�\��/�7�G��~sQ�S0 ���J���LM7�3�؞�$Q�c-lg�X�6$�h1���̒���5�W�g��8�as)��qG@Z��4c<'X��ԇ�x�v'���_�� 5Pv7���j�����~�.�1�����&��U�ҜQ�.��Gsf%p�@�o����O�x���Կg�<�tܵ�9�~r�e��2ʬ>Vqo�""����C���Y���E���l �>�������&	E�zu��!�r����n,>��9c��?;3A
�K�o�]ىI�{�g(y-��B�\a󖻆�����h��݉}�z�q�%��3eՁdZ��o;q�ś�74ʛr�I����K+ܸFj ��37n���OM9E�>���?%�k ��.&�2	�B�����(I�BX^9���Տ]U����V���R��o���n��"oj�ŧ�mx�8�t�W>̵�
�1@X�i�1���s���eZ,����{3*��N]|WĴ�cG�M]�&D"Y�[Z�]�%30�K�U{��n-�i���Na<]DI��)���B�޺��1�xz�W��{���k�X�M�\�Y�[�e���Կ:��1ʮ��Cq�-mð?b)*,�}�|�~N�cz��kb��NP*;ӌ�4j��-\Z��X�P��m�� 2&��*�Yߗ�Г�1��m�k�C�^�|����Y7�]R�0!�����3!��2��PD���rs���V�¾f�i�;�>��@#W�3��TU�I{�̆���:U�mi��;JB�`�.i-�sf7E͓`-��\�MnU��J�Щ(M��GV��ۈ�R�M�Tj\��� ���7��kƬ��!@4��ޢ��QM_�tK�"SX���U�I�h���%�G��;CU|d[6T%�͗0X�;b'�1���s��i�඙±M�D�Unj7��_Y�s�0E��;$��1��÷h���ǽa��=R���e�\C�밚 �����h�R�k�?q�:��KT��q�ʂT�0da��P
�H��(ZL4xe�g]��j�|����麁�L���;��s����i(�=�j-P'�Pi�#1:�B��+�Ƌ.�qgU��� 7���RH$�w����L~�Q#� f�V�!Ƨ��O�ĭD�I��F+L5�q �:�p�H�j2G�p���k�4���b�\���
BbA>����T�FN�~��0�͖�vB��dXp!r�3��F[4ߌ��]���@� y�"ճ1A��vY�ؔBi m|����� ��S��c\ [��5H��ͣavkS�C�ud9�;�,^�:����?ʆp�!���%�{j/���dSs�nA���|����+��'�)�<� C��d($����#܃�M�\���$��_�jC
_��sƘm��ԇ�K�%呤�?�g��kWd���d>~�-w��c�Ac'z�O�����G3��'o�ŏv��2��c�xb�yN�p���eS�D��UFQ�4�h�$�&^�/ݚ�%�%\:d�wn�{�Ɵ1P����*hڢMsUr-��U+=���V�_*�P����ڠU��p(2Z1D`�u�gȲ��0P,���TB��S�L����`��E�S�θ�R��nK�8�=K���g;�ǵ�tj��Bvv���7�<l�����g ��RN��; )�9��ȆIT$6u��ո�&�0����O�z"��{ <��㹦�8���O����3�(���K[Z�9�"�/�u����޴`�O���l2#a��K=�:IK	�g���s�������E$B�ʀc2�k&,��Hu]��6��H=��o׵F�5�(˂T����W~~e����/T|�2��5���:W�[o�����^%_�A^�_G�����Im�`�݇j�9Yl�t=����C�<P�m�6�P�<hF]+�̕�R�_��M�X_���B���ū^bb�4l��x)>zi�w���E��+	�.�+,^�U��������4V�F�n��ofE��P�I9fa�O4�y���FĠL5�z��G@��e�(�f�lXüEGf9Q�d�Y ���Z�}�4�����M���o���j�������:b�2��UIx�N��3�6Q�� �{ƻ9Ya��D�g�s�R�rg��0r�
G-갮K n`]�B���	��T�^rU�u�Z։V6��-Z!$M˅���!">���>�#�w�r�z�>��ٗB'ZeX�v�E��2i�iQ����Fd������RN}�n����Nfn��J۫�_b��>!�y;� f�re�����,������R��a�0:����$�~��L����ʂs6N����]����g��'��>�k�v	 g��	k��ZC@���*i��O:�������x��vH��0���h����pD�]/�濔����gBd?xx���j�?c|Ӫ���.֟��s�X^�(�I��������i7 �p����0��:�J� ���7TPdR��A�6��.a��AE��L��F���s���A�⡸��J�nq�is/T���D��RV��c_~�G����F/��7�l!�R`M�gl����qR+$�*c���X���1�	vKj#���*ccIk�߃|����ki�{��v�WY�ę
�T�Nb��9p�4�m*ˑ7�İS�dG_W5}�&��2�z����;U�D��g�S�ԗĎ  L�=�+N�!y$��/�E1�<��
B����I���E���2���L�ٌBE���$@��>�q+q��7G#;i<��T��D9Z�I���	�%�~���T�'䨍T�Q���L� ����uM�y� ���	�^��0z�wBs>D�W]�GV��$T�+��j�RI\v,�)c;C�_L�������+�߶"cU����rk�;�<�I������&Ơ�����+��ZM�h�;j�pF�|�MK!d@�-�Ƞ��:0�5�R̼|I�"�$�Ǒ��SK/y~.�t^�|Z�����2-3~��b��2?g-oM G3���s�%�6E?FVI��m{cM�����ʇ��\70��i�h����*���lKe���#�_ Z֔�}۬TO��NH ޽K�S����v���>�_���"UW�Ӄ����ZA��2�����vgp.��R�;ؐߘ��p,���Dۚ�Q�S����òbN�X�]�8�'��p5g���9�RB��|X �Kح�i�V�!&W�����~h��t.�K�)P~;�������C�Np��@�/�t��6r��c�y?�'�GhG&zz�ښ�����	�ڇ�4��Ts�>��q���m���M<`|����� r�^�O����f�fai��^��0_�/��F��}~=[�͉��S�J��gE
	����F�r��1���'�1���LZ�Ѭ�ퟌH���c^i�}˟��h�0��V�Y�G&�h��3U21��m�P���.c��RwRL��"Q��goM3E� ��+��0�a)�Ae�GJJ����ߌ�ӻY�b��&��%Q"���/���6�{I2]�8�����u�j���P���Ǻ��o�P�!!c����07cfqQg4r�Ղ��z��#:Ќ_��}�چX?�m�H��%�l�e�^3�sHqTz��=��/�K�/���1`F��7�d�(҅�$�6V�>f��$u��y/DX�����)�c�pĺ��%�h���8����GP0��y<��E�~����������ѷ�e�fzy���r��Z�.�b�jjvK�;Ji��Y=�ݖ�|b�j#��E���"����b-ε>�8��9j2ų^�}T���0�V�=mtA>��2D	�}�t6ՃQ
��G�]�'�TwL4a�w�-�D�M�Չ�ȝ�k&7S�f�w�"�2�/����1A!���^ޔ��cr�K��k�����Y�^�PR�Ii���Έ�
�絵��C���?ec�Aca����ODq�ѥʈ��V��K�u�y��~�Z;իM^q�GT��O"QJN��u7O��d�U��`���S`�b	U�_/K��~�􆀽�D��o�n��\
mz%���M�x;�_Ж��8y�bE3N4_(��fuQQ_����|Ee����'�ϒL?(E���>s�jxAǘ�ه��v��Ã��K=������6Gb@P�4���?y&*�Hv9����u}ʐ��he%�lgb�tp.���\�y���g���l�l?�@ɨu��!��nc��T��� �{�W�2~��t�^� �C�9����h1�aw�Un�O:`�q�m�Vy���E���]�Ϥ&���������	�6����k�|��o�h�#�b]�Ni�"��͕3px���������A\��tx���12�(�0U]��� �pF�v |����(G��)k翉���:Z�^?����w~/�xAC�*'Z	?V4��o&qs����a�����Q����q�jp���3��{5UU�d�<Աì+�a	����Nv������/��&Ȓ�N�K��ܤٟR�� �R�h�ډ��%�:�y����oKq�GE��ȂFUH�	s��Z������������͛��	^�m]0�;;fǎ�}($�"��#��\f�KUʂI>�al��S\Lٜ$3��߶�Jc�*F�c|,��l	;�ʋg�՘i���/r�o��܉���ƃ+dw �#��r���ŵ�,�vuW�nx%��l#��L?�a���\�.s��F�^l�Z.O+����frE�1�L'���T�D�b�Y'�r`��ybc[AM1�#5[���A�49�gyR��.�7�G«�>[4���c�P����|h��P��)�����6Yl�K��� d�4�"BCb0+��4����uj_u�lU�R%u��:锊�9er����c�ȼݻٸp��Gt|t5ɨu�Иx�����C8��S�*�giIwA�l�I:;����1C�Ł�FS��m�F6��&}�������׭���]�U��]������^%2���5{qI1j��ǽO�������,�ҿ���DutT/`}�D�I�śFo��ꓯ�� ���On#���W=	\�Jc��r�KpD��m�u�.;̇܄k�~&*f���;rLw*ïm"�w$;(�mzO�(���"W��>`�JW'c�o]���Л�6~՗!R�6�<���?IG7�KJQ��<y|*/���,t���zÊ�F��V����ju�	vҪ�o��8�Z��V#5�T1qP�b�Y�j��� &��W���qIi^��)<����p*G㟌k��0����N��( A[{C�s1E/΅Ǫ�c�C�
CV���W-�k��re���1�հ�@J���Mq" � ��Ȫ����Q�Q�}�.��4�
�Dz�\m �AE����b���K��Q���doEb��80��֎���ﾇ(i��"_�F�����q0���u���5� �����G�V5��w�U�U�L�[�q���B��c�ȴyF+$Q���-d���
W	��&ɚ�'�D���-�u����	 !��G�l��y6�z���}�C�q<�� �0�m�z��;��[�ȤY��)�>���}'����+H���	�Y������J₷�AnshuJ�w�y����:�+�}���(Q� ���If�\����;	�ױ�cY0T�� 'ֶ	n���6ፔ���#|���JB38�����]i��� ��z<��F��%#В�1W�9��.\�g�*>TI@�ޝ3(��$���C�zq�7�E�e�U��Dɗs~�Y]3�Q�N�^���v<(؁�@�"��AVT�����%�vv�6�<qH�c�sb������Y�`��%�l���1��	V������31I&�-���S=XV�R�$��Y��͐M��_�~s,l���&�⣇p/�N�G��݊?���1��؇�@�n?����GWȞ�2D6�� o���4�`�'s@��lj�i8���y�+��H�{b�,�%�Y`����B�4@�nd�1���
�%�B��*��Eۋ�P���Bb�G�̰��������H��īܠE�\z��d{J���,Z��AD�ڹ tJ)�E�:k	��W��րC�ڙ���O�6#15Y;�T�[u=+$��=���}�ߠW&�Ѱ�L�����ks�ۈ��aJ����e36�,PK��/[+��$�؞	�_��+��!v����H�	�vJx7�iD�z�Ld�K��7��t�pE�A�qx�|F�2�܃���I�U�	�	���K��p]�w��ԊtA�Գ�A ��b�����7��#�{ws�mK(������v��·�ON![��9򜇮	�G�=�T�����-���<����D����}/���4��V8���]�֑�L �+�&�!��E�J��Ι���%\�;��2Eט���{e�|����-vgƌ8#X�&[���ެ���Z���+ȃm���3UO����:5�w4��uҁYH��c�a��SV��-b���]�d� �.�>ƹ4�Q$1{�2��?S⦳3j[OL�(��.�}Jj�x�Ө:��E� ZɃlt�������}Z�լ�*;b�]T�k��QM�����>���IQ�+ ��vs�����yy��:�d��EH�=�<g���Q���K��R���Ռ�/D�'iQC����L�l��&�te�81�$���o&x�J�:��	�&�������"�h9ވ�K���Z�C�m`bd*���ֈ.�:�8OK#�N�COO�3-�Y� ��֘���;�_�w�}����f,G7\@�㟨��"ۅi��`
��a�W\	 X9�iM�;�y��>���<Z��h&�>~� Y�����=
[�w*�(�CI��@�j�d��
�r��� �7s�08��O��N}E�Z;>��TtWrBv@%:�@��$	�1):/MqtbN���������ƭX9� ���=�2~�XI<�"�&_�Uޜ�<�ʥ%�Q���֙~�y�r���U������f�����n�\UC�x2k��\5����:r�w2|�KJ�pe�gm�����PZ��m�Q�¼�
�{��a��q]��� �%vS������õ^j�X<5�̮rs<�I�\d�6���nV'��m��Gih��;Q�*J���.5ŹTs��_R6]�!����.!��h��!sf��kb��r��f��0!sҽlfzJ`�f��D/2c�5�7�+�g)�N���Bo�X��ס|�$��v9n�J
���
�7��Z�oS�������?[��'
�Oi��6�T���f���������._0�1-�#��M�xx3,�LVf�M�ؼQ�%X�;!T�t���Uݵ�ex���z��K�D���<u'ws�8r����u��X�g�L�G��qWA!8��a�@�~�ω̸�x=��`�U�������d�@���7�y��u/s�l"��b�W���L����ĭ����;sG�*�V�!��z���d�E`�Q���򩪈�!�9���o^�n DZ+զE�7B[�3�;��hd�NȎR�[ǰ�j�!��d��!t�����3�� �;p���~������;%�OAa��ϗ�Cx�F<�;��堞@�!kG{srQ�����5���H���?D�C�ļl͊��3���K6��F��I��ȑ�@Kg�^���^�|<+�!D=9�7�È�t����2a�
5˚w����`�_�ݏ��F�0�]�x�ŗ� d8���&����~��6���gl1��b=���v~ 1�̌����X� ��X��G��&چ`(��)���v!8�9��Ơ4��I�CD<%}��	K�k����P}gԽr2`�Bs�&v��V<��v\Lϯ��zs�l���
Tjį�R�p�&Z3�n"��I�a��=��Z��bp�W{B~��	�BBg3*U���D5ᒯ4��e�[2a8�X�
0)��R������c̲[[��)�39�f�����Z����� ����A��^��`#'$�џ�f���hVx� � �(=�?��	.���K�_���6�M��N���©�6�S�J�j����W:0��#��n��o
�V͠����t&Q����5.�"fX��xZ�\�bG�L���o�.E	R ���1W�#��u��:<�r˟Na�PJ��wPI�< o���%���tW 0ޥ�I�K���H��[')���>��"P�d~w��Y�P@7}��x�Z��м���A;0�����ܥXQn>�+X�i/�/0O\�C�2��UR�_�
I6\L	Af���� Y?#����Y�{	đpF�pO K�aڹC��ϭ�HKg�K���ѓ!��wN�(�_���!��3Jȸ!�A���G0��Y�}& -:0�J�K��jHx+_|w��k[z�(ˢŠ�Rr<Un��߬o/��#4w���b��d9/f���<oAl�F�SX���:`G��-�Sln���e	��i'�ϾX.�)g���y4�確��-r�+��lU=�p�(�Q3'v����SL���R>B���t�&<`��E�eC���К�K��T����ti��y"��@���^�c��d�ؕ�&�D�~Tw!^[uG�Sj�8^��j�QR�f���0(z�9�iuQ�E��w�r��a�.,_��h����D����������ޅȑ�O]pCs//A
9�K�D͗;���X��/f�g���a���.�p�A�-���^-V@R�z(��F�?�KA(���������<�/'3���� #BWfm�E���%E�a��X숖�C�{�2��r�?�ȑB骙�q�я|4	D�q��8�\Hu74��d�Ij]� ��S�?�m��`�UJ�]���+���G� OV�����w܃d��f_~����|[a�/��_7�:��xA(k8�:p��*�t��F�������vSK~`��H��@v@r�8|&�y��8P�{��F���7�4��ފ.#�L\�X�6�UvW�pg~VPH�:�	��#7$t���4�|\�;��&��3�]���3��Z�p��'�1�l'�U����ʨ!�Ws�y�R�$<G!���ȳ2P�%+Δ�'��ŢY-�����h:`�i8�xI�R�:қ�t���xb��q���Du�|k��K$��+(.9gK�fNe��L}<{D.`T��Jij���d8�7�D+�9�u��i��� }�}�k{]JHyk*���.�d���J��Ǽ�:व�ݠ�zu��f!~NWg���#�nM{
;�mz��k������,�`ŵ}���;a� m*�B��Ţ2�3K�����F�!:x��Y��r��)�c%� ܞ	&g���
9�..��oo�6 �yK~3>k��o��A���̿�Yug(����Y��Y������*V��.s��12ԓ�r��3+7�����A��ǓW5�)��)O��B��p,�jnE>a�Yl��o1�̓] �Ѝ|=3~n�vq6�$��~��h5�*q�ͩ+�f�Jz�N������}+������U���q��h�N�vaA��c�����/�o{�� V��*i������P?�1�������b~g�M�f\���-0�r�
�w&^w��Η�q!������_�\!�Zi�׶_	���e�W�N�� M��\�W$����|�yH�#cϞ���e=J�<�	is��.0�S�C�0'p�.P5�!� �-�7H{��;�L'$&�G��Z�I_{�Q9ʦ[��J����D���,���4�F�a�0jgЍj��ҝ��@�)暼K] �I�m/.���J���1���_-�Y�SO��i�[45����F9X[�\�~�聕��ٹ!�jvNE������� AU��y��}m����G�����('9n�nz�m����#̐T��Q�'�0X)������wJB7���43�N�"�o�b���r-�4��F0�rs�S�r�â�q���)�izYj8�h�-e�d���7Q����O�0�K����'�̡�s�;��fDbU�'��ƚU���7��6����TfkR����W�X�#eSJ���q	2��k�Z߹h�K)����Z��b��ѢR���Ș��p�r�*
�����UdR�����e�X�7������T+%��,T�IΗ�i���������)a-[��E$�
ǣ~I��o���U~f�����(�:�ߌk_�n�,�6�LЃ� ���W�/ő\t�P!RP���X3 ��ҿo�
KOR����C^\���~���fa�+���z�>�H}���&g�\��b�b}���jJ�m
�FNK�x�4�fb��5����6Ο}���F
� ��+���䬖���.�b�����sі� J������ϒ�^�L���G�r������C�#�E�k �:�q�x��k�tE�	�^S�Ȳ�] B��+!r!���P��r��/=��F]9zW�"��><-�{*�$H�g��m�\e�D�9��U���*��ߞ�[h��(!����|��P�ؾ"b����I`�v����q������3�.�Q:��6��@��S�'4�\��8Z8��#ML����������o;e�N��h��q���I�gPb�ޞ0O����=�~�<֞P�p_4���ذ/me�ŗc�m�ӪZx�+�1{�#�3V�)�|2�UE�����HtIz��\p�h�w���Yk41�M*�@�o&9�4�e;���,l�2xS�A?I?,_��u�Lr��ޅ'O�Ap�\���ڳN&��s��J.�#}�D9�:r�F��&�-Q�Lw��U���G����}�<��6�y��$�Ua�N$�!ԏ�Jsora�-B>)4�pݾj���$c~�Xx�- �o���h)����2��|Q��9y@�9P45t��Y���� *�jsu���Ps˻	�+L�q�OB#hZr(T��Ua�'��E���]�P�a���~L=����[�S�o,4a��J�������Lh�I3TmT��_��~��#FϷ4m}��;·��I�ȏ�C�Z�B����,�N�y����=RT�y���;Ķ����_&��)���J���M����#W��/h���;R.�����#5,�����a�^���͐B.�i�W����%i�v`�!-�f6Ю��FcG�S���'ר7���5���g�*�S��|�Y��!Oz̴1�c,�bզ9��qV�Tg��������Ys��<>��V$�
\���%P'�=w9ڀp��AӞ_�v�d*ί�{��Id<���'��¬k"�ݳe�v�R3��HN��4�Ü��/�DT~�9��(uMuF�ѵ3���ͅǥsr��Q�(���$m�,H��<���N�8|�Ms0��v雹C�Ñ0� ��������1��'�*��E��g����\���]���j����ؤ\��αc�p\+���%���WJ�� G۝7T�(���6{X?:�˰c��2��ǃ��u~ӕ�c�%����)$�2|9��"�8&Eq5(�fNq�EJ�orf�����~qҽ5��y�h����'4SR+o��{�+�>'����33V`2"���	�ҽX�=�]z[`7H?�@�{抅�p�Cq(�\����ɳi���/=��W����)Oo�z��X���`5L��yE�=_ 2��Ɉ!�˕yJDuPf �@Q�L4�d�u�-E�g�9* e�g�p|&�a�&�0��a�RiȭL�������}�3.�,�Jr�~D:�DvT���<�<%�|R�]��]Ɗ�P+�8�Ԕq��QXl���K�6���h#�y�<��K��Q�X��ux�j|4kX�HN]�D�ƬH��g%`0IA�~�Ų
��Ĥ�$�G�K5��/wR
6��4&�>@Y�2�ܥL�o�e��A:���@�ső;�JFr��Q}�8�QBy�v�V6����a��gd��S-�]\U�Yp��0����T���eHh�֜�#Tjp��J��x�@�X~Q_gF�t�v}q'o�bOwQ�����}��O�ν;��E�U�6Fu�esF\2�^PR�H�q��]B��O���M�Jv�Q��A�|��.,�!���I�m�r>�fx$���� $]"�F턬�o�R�'�1�@ �'��ςƟ/d�����]�F�x��A�|Ԇ�p�$zV�y#����`���j���du���ŏ��匞��0Ǔ�r���(�G��{��b�B�'>]��d �����D}���d�0azn�j��K<S3yΠ�����S�<�,H�$�#��t�j>S�x��8���;aM��L�I�ӷ8� �li�]��v��}�9ݿ�12Ec�oHk���E®�󝅋t4( t/սΣI�=%��#A�������y��7'��x�����oE|�Q��L9�z5+�I���V�������̯���#�K�G�^�X�0���P�Q�&�&�T!M�L�P����  �`9���ԛ�#�+��h$�����3���e
�N�M�n1V,�"s�)joM�o4{x�2I�+;���S%G{��R��{��N@�Ҥp/�D4�u}lFն�p^ƿ��Q�9�19��&�9�X)�]��R5m?|���ALJ�K��=��d�TtЍ�`ʑ�E��t� �<��e'�n��^FM��r�&T��t�4t��U[	M��%��V��ucS٤V�,^�}���(?�n�9mįQ���W�� �s4��0\y��p{�U�9��L/:t��ϝ-X�?��O8�G*�q&:�/��&����)��o������m��$8{ [��4)"ʝW@���{l�������Q����"�n������|�ok�D�RQ�������̰ e-0/����������dڼ+�z�t0] 2�����0��@�u�;I�!m�nvaC�z�oC�G��A��H�F�0���x�ԇ�^�\���zT%4|(EI��"!͹�Q`
�xV(ʉ�1���Mn�8��&N5�{w��{�g�08=i��3RJw(P�̙>)��][�I�H��e_s~,�8���zs�Xh�����p7�������zL����Z6��DI�i���x�Ǭ���8�V��(�T�}��-���tm(H�B��Xb����hR�B��v��"-C��X��������<Ey��V�3�PB�J����t����~�9z��}�l��祐E�P��h�E�H'���X��W;��lQ���q�07w-Z�X�*����Կ��
��)��
x�M��jh�ͰiH�x_	U�>(�4�B�uRW7vkTW��]�,Xr�M֐җ�V��b�2����>�l~$m�-��៪�n��M�T�Ҹ�
��
. `M��SD}&��s��}k_"�׋s��!`�7T�7�<iS��x�Aߚ� ����|`��%:�:�Y|�	N��d,z�H��\��O�/�g�)���	�FM�s�z.�PNc�5:�y���В����_��C�
D�üFK�D\3B���������i�`u��`x��%�4��m����d��X�����"���J{"�I�A�P�jB�=��iT�9"�E���~(:����E�B��u���G��V����J����`�v���A~��w=���ʂ�r�!H�qO*�bda���?��<��6��2\!-F���.��{�J�n��Ed����R�70�;z�����
=/ h ������y���n؄�	.��?�M�{C[&�y
��j��*8�zUG�'�Tv�,Q�uY��7�l#0qb��4�Ķ������J�<d:8$[I}r?Ԝ�c�TB�M�H��!:�B;�~��;Kr�@:�#|���HG;I��/ ̹��+�g*�tD*bD:d�����"�;�	"2s)�ѱ�^�Z,�'̾Yk�|�n`?�rP))�"i*:3�H�m��v����RQ� G�m@�c�M����&�8�󤺳P"/��7�g���m`\����_OVΩ���ݎ�tH��x�?��م>F�CHE�(5�v�1�&�'�~[����T�A6=�5���*t��\�ےvB鴣���|Fga�>��vYl��-�0��1I��r��5�E%Gl�Ĥ�V�\�p�1؀�U�l%���4��C��ܵ>X����#a3���X)J;
���)�㊌�ȸ�0���o�N�Ih�I������"fa�����a�݄60%��}�ང�����^��4��KR|�HT�~��?+>���L��sg��GME/��	��J7k9R�2LI�,�I��LY(n��}}���d�!��t�X����1
#���Տ]�]��U��v�����ci\o8)�2:ܺ��c�L��,m�IQ?]�*�3�?�22��"�\[M�v;q���>ɐ}�ԍ��?7�=1�8\�
̪*LZ� �&������7�N^�яq��r#H��.�-�����`��7@˽�6)?���g�.��ܮ�P�u�=)~V�R$����-=�;���N��zʾ���	��wxl$��(Rs<�Cg?U��Ϥp���^�vr��1	�n�*g�|����[Dh�C60r�ғ����Ո`V��?�+��D��;Q�YB�i���
��o�9U<~�����}
ߧ�V�6����u� �.:��wI�����b��2���H��&��-_��O(2<���E�������yUB�壦2���6)e�:��pkX��I^�����N���K�r��Hȍ����,5�(/�9����G�`OSq���/���-#r�ER���}4��M��쟗��<X�>���Lu���.�/ጸz�dᬽL���zU ��l�6XG�U�S$��g�}�Xx���v�p�w��n�]"S\�h[�l��
��g�� ?�<��)�"�(��)3d3�+������Cl��@��J�̍�`�
Eu佱@@ꈮ�����m�	,�H[��Ee'����1l��<���h�\�p��JG���Q^7���*~a����6l�����D��t��%Պ%Ĳs���7��`�#�O�?F��9~��/=���Z-;R�H�OЃ���9�O��m�ՉQ�	��^�F�E��@�޻��pXa��8�s���h���|��W�E�x��lq�!����S7ȍs2Gn H]>�[ 4���گ���EPj���Q����`�m��o(��!��7�3�WD,���29��͈�Y�$� Z(�	�)��BϹ�FOo5��^8��K<(azp�$̩�*C!l�֎T��O!/ɯ�X�d�W�Fm4uiǿ��L��{�z��!G�k)ݘm�)1r�Ll����<u�Q�>���g�J�qܺw8��x5��s]zD������B�TaJ�����$&�_�h{�O�������Ȑ�:���b�JH�
��F���J����Ė�>�\Hx���
/i�4�G�����	Q%���G}�_&�o����b3�`���Q���E��oGU�M��$�z]ڡCV�����$8W@�o���:hf9})���d�?���T-�5�Ċ�=ԝ>�nx#y�7�3/7�����k�������CG��E3�T�@�e�lǪ����A�O�XY�*�pv�tǱ�D�*s0��Y��5p�f�E���1������D��_�&,S殗T��Q�.����D4݈�5x�[�ݹ�I��[꟬�����C�Gk|Q�i�j�5��X ;d�e�'=�zo��d�f�.7B�M��
o�hK�Yk�h���Rn�s�I����sJɵ��#Ƌo��a!Z#*��5�����#.k�{�9�v�N�`�8.���%���5i�a�F�	6�<�v���膈�k�4Z�s���m8����Ȓ�2��h�ɻ���ӌ/` ��f>�`WI�lT�&$�N���\�C-b���m���2y��zZr��׺c���C��L�HN ��o�|�_
[��HB}`�Q��_�ԋ���"�f!�B�/�� ��W�S�@��q��=}��1K��`~�;D���YZ\��=���Cd`&�Q����<ZIr��
�I���7����8��ǳ�-/�EJ�{�,1�J&�5���=�m-v�@=���$�|!�6�lҥ6��֮/G֞٬6c{��?�����4��
��Rbs��X��圚�&�ZpПۣse��S�]����^@�s���s@�\��n�,�Zi�k�-e��?ˇ:ɞ�~�M1��0kb��A��@v�����t�~����@����Ίf&��؅�1�ϡCڹ+�|��B7[�-���=��^vա��S�ZLk���/̗!=��
%����Q�WSI�Ĥ>�V�Oy�7Ƨ���5����	�n�m��^gP���3q�r�[����RWd��X���0H��[Ļo0�L9m�N��1Ǡ��������&�hऺ��}�cj!c2=c��W1�{�Fp��s��I���<*~�S��
�$�g�ڐ?9��Ą��u�*��H��5���ņ;�Sa��ͯ��§� ��e2�j�2�x��_Ԅ޲��An��xn�ƾ+�mB���}�_���J7pv��9��c8�C��b\����^w`ͪ��Dῇ8&^�e���� �i�S�h9�x���5K�mk]y>c����t��<U�edl�8�yI-�U��Jwvb	���Id~���?�Z���8+�3x]��L,h	� ��x3��^�eݼ�M@-"G����&��G��&����XVs�{�N�KYw�#��u���,��i��OQ��6K�����2Ǣ}�v���5AA+��^W�ğh�1�����KD��3m���Kw��a&~��'�":]+�k���)�.5A����H��'ͯM
��=Ny�m�
�E���ȭ�Yt�H>��]�	S�f�q[V'K%�k��M�mne6�Ky1fw��tb,��6��>�je�)�+��T(PS�?��*T3��pZ���<�%�x�?f�A|w�dy��o��{kO���	��+"k��/���2N���o�<���Gm쉷؋�"C��L+|�rǵ�MH��d���*aW����=N-��π�Ґ)����Z�Ռ���ll�E���IsI`U=��4W5o"X�e�q��T:3�a�i}�d�����oz&o�
/�D���c������φ����~SL�ݽ�wR�.�����u���}�Ԝu%��Qa������
I��c��Y��L�������s1��v-"����)�q�+d��,�uQ�E���|9'��p���x7JȤ��/��Jz��M(ݕ^t�Uɬ��>`PK���_̔�_JA��l)>D ��O/��΃�WZ�u�|��JD,�O��Z\��n�_h�.��(���W4��_M{�Gaﭷe^�q�F��X\�KF>��<��a��Y<�T�A�؁;�y��h�F���1�E��RQ����r�E��k]��d�RO#�0R)�G��1� [0� �m�-gsP=�{Mht`8�w�����k��NQRڸF��uM���
,+�����3v�ig�fG�����{ӏ'��&|ٙ��ǰ6O�^��c�$�4� Λm�����ub4A���1tܫ��b��Q�> �A%�4��E|�Dq�R�8�t�H �e��������M_}�bΖ#!��g�E7#U�q������	�%<n􁌳$�H�6�ߐaew����@ajw�|޻���Op����rDʍ���ۘ]�^zƑ��`�w�%���Xd�˒�+U5}�������hPr�di��s��mt5�_���֞���۪Db�������B�]�P�,��c�D�޺j�?�%̱e�s�Ʃ_#9� k�����k�:)(8�	��. K���Ǝ������P��M��:s�j0�h���-k�oպV}�E@&�
M&��iv���&VH;P=�@4@ ��/��u�1!�*Xڬ��%��f�pWMĨ��B�#�@
��,����}���u�T��G���+,�G�[L���)<�</�0��Ö2�+BB���cԥ� w�X�l�Ƽ�n�9�@,b0�c�����A �i��C/�n��[�'p����￨mO�Ol?�@Wg�il����W�<�4��۲�ycQ4��"9����-�� ����/��~�#0�eȒv�Ze�;&�-cn�a��Y-%��y�6���\��
�]_NkWs�!U�72M��$�'}f�ê3��>�&�Iz_����M�G�ݝ�頛� �l-լ�r���j�D Xukw�ڙ?'�ȴ�Z��%٦�ث���ls[�n�8�B@`��}�$a:~���*4/b�������_���t�$�oth#HG���$��.�����q�u�k�_��k���m�z�t��B��ȧ�ٯn���� 4�;���音e��q����rݐ�Ϛ�SŒ,rX=W�/�?�I�1�bj)ƽ���I5�D�Q�|脛�)�i����V����s��Ѹ��(�'n�J*��o�.�B*&0E1��M�w�c����'��dӗ�쵋���e��� ���e|���*���~7��#���K@�O|a���?KW�4v�bV�v�i���V��u��E���Ky[���U0�C�4����A�o�]�m,H������@>�<��Z�����2Q�G��v�]��cCW絧�%Y�h;��w���M�G 0�)�L6{Z��u9��?!R֮i���ķ�(���p��2yx����'����
~x[}��ʝ��x����z��@t��s�w��9 ��-�~�{��=e�����SEl��c��bi[�	�^5��s�&�{[�U�0.�d�h�bn�L�Xe�X���sY����w�fGҲ�lI%�4���̡~+Ezȶ~/��A6����V��C�k���y����}����&Y���O2����q�n��%��'*Mʛ��O�]yT�_Sû���'�
�K��џׅ�:�䰇{~%���*�\��B,4��쮬Zg݄B].�y�;�kg�䜛O�Ix���B(��'G�d�<�,�Y=���J��J?_ �7�w��Ä��4&��/��3
"v+'����恵����W4��E�	$	=|�~ߞt9�23�aD�6���5q�s���o�0�|� M5�D6BE�`���OdC���1�U*�w^�qM�R�}e�,����
Jd�O|Q��c�_�����X���eoEh�����
�[�
^uT���8�ﾵ?��i�/Sȡ)�3���f̳]w6�j��b:��V�(I��7z��L����P
�6}�0��9u�+|_���9X[̆ˑ�8��{�8j�L���`�b/0p5%�O2ŵ��[�˾$1XmR�jl�)���^V��39I������^c�.�FD��k�aV\���nA+�Bg�W����h]����Dݷ<!�P��/b����7:�ۜj�&!�¯KǊ���.�]�M���N�z-?��ٰ�)�x �{K���
/e�e�D�y�s>Ȃ�
u$��h������L��ʠ4�`lp-&n�6�H��y��_%��� �S���E��F+dP>�^�+�a�1��h��T���\ް��.�(7=EuJ�M7���*?�K6���5F)f2_D�+X��K�,ݼu�7���*W�?��2c'��)������=2,�������Te������P��ɑl�4p��[p�d���+{�����KA�j����~G1�i%�h����G�E�t��&���F������Ώ1��.J�p�N+2ud�$z�s
�!�k�e`����Z�s�Y�9K"�����b\���%���ցؤ��d'��+O���X�R
S�W@D�i���v��A߃��\w�Y��X��q�}8�C5P֛g�Υ�ח�l�z�!)��3��ր� ��eó�:��.I�0�G�O~5���p�޳
��s����0.��	�{1�H
��17vK�i�� ��J���14�KT&w�%P���e'Uq�1�.%���ko9N;���������|��&�ǈ���/�Mz��ٞιE��9��@���xhwz��f�/�����D�0��z��������������%LcD4s�䩄�����WZ�?8��|�u��W'g����+�dWǐ��w
��g����06-���X����u�˲x{��|�9rG�]k��df�y4�팥�,ʺM�3�XV�"P��-|�P��H{�
�
�n�����u��p)���K�Ү���)��#��6��X���G>��3�i �g�~Kr�c�wW�o�\f�
�{a
75����D�/�_n�׌
H����Z�����e��N�]ŀ�g�ڋ$K��[�m���f{o�gqB��D�T3#��웎r֬Ju�S'.>s��:=��&�x���Qi��O��Ŗ+�TBv�"��I�	|0����x s�u�i1�e���� C/
���$H��֭�������m���B�*��=a?�������D䏋��d�)���!�M�(�����C��jjx-���M��E}@��4ZY�<��*<6J���� 1�Ol�ٶ�0RG~��E�8��S�?���4�yf�I�"�2M�2�����x�]�gry2�e��Vu������}��%�>�	�H`j��K�F�!U����Y�ߘ��0�W{�*lˌ��r����]�&�Xy�<
�;M�|��?]��|`�>�=3~����,����Y5�_�`]�|Ӥ��>%~�=OM������y<��+��q�� �Z�<lt��׎���vq����4��2&z�$$ r��Jgp�=����2�Q���(yw#�c��PG��?�
Go��"��s7�D�8@��5�	��1^����R��^�����αg�,�`�����(��9��D��dbM"����x�&������-}��:�,��EIG�_+NLA�!L�
]a�6 ��W��
���9��}���Z\ǘ]̹���e�������ې.��<)���V�V�����)KZ�$��Pg:���9O��:�����S�-us�W�.Яy�-_��#�N�������2K>i�e/wB5�v�����G�a��Cؼ(um���?U�נ�^��r�d�����љmWo�Zm�.5"�z1wcU��P�������ij꿳2G�-?[�#�G����MO���V�^]ج�=�*k=�:�]v�5��UЧ����:Df4?��c�=_\�br��[�X�v���f0��S>z�_߅�*��O��]w=�u&(M��6o-�VQ��O�,iԅ[������~�?��8ǖ ��2@'�P0�#�T!��]O�B�/(�?�Tn@�ʠ[$Wс /��n�mL"򒂗F��mR=��<��Y�Ħ�1���89q����QB�Iq��~Xr�N�m�}mC6q��>���YN��DJ�e����΄�Н�A�ˆ8Uz!�Ky��&nca����r���Hb��Sq��#^�.D���6p/6��t'+i��Z2꨺�Hs�����R�`�]��`m0��Dt���ޥE B9"��uИc���)��PM�ܽ�u�X	J�I~�텒���?>��:}��Y��}]5����+ny�Ky�KLh�ሃ��Fg�Uk������p.����R��#�����Z�*H�
�5���s���A���i�D�%���K��9�gc���B�f͸�6M=|#�ÿ5'�
-[�6�����UȂ�s�4�<A��Ex�/�>�+�:q���Ѿ���si-�Ϟ!�,�1}1��L��������DW���^� N�ƿd���c�B���ﱕ4���K�O	R�2�>ȁQ��vRȸϢ|�4�&��'���Տv�|Z��V<Mt�D��k��c|�X2�jP���Q�	�IL�\�R4�V��Ϧ�Ș��x��2I#~���ˁK�8s�bꏘ��	�%�q�Q?����N~�p��,v�+��g�Ѱ�=	�n�n�G��Dr�'�q��.�	`+��+[�\�ҀhG떘��m�>�4��!&�&���vx���S���W:�}e��ᆭ#���=���|�qo]��2^k�u/C�48.���P��ϴ���8C��9�Ϲ]��'�n���~G���A:�@�S���xӃ6�FvFt���R}�����
j���ԭ�~��oM�ěg��v��w��H�Ϩ-�����u�(���-�u��E����ʄ�"��� ���wrG"/2������=Z���|/o�-%uCӞ�[��
JR� !����(�˕���uk�@lbld^��/37���[X��OW� �7�{��OtT��]��ٞq��4r�&�ܜor��Yo��~���Bw�|7���ܫ��,�j�M�g�O��|�"ևx�6�u��[>���
@`�Z+-8�c�'b:��u�a�w� ˔�����>y� ґ@����猷���׫���FP��Y��-��]�rLt\#F��\V�NG������4J�_�#e�1��}���<m��W�²i��_��?my���#�\+r��8�J�y���7`&�y���טHxh�Ո�v6*oI A�����|-��in�����m��ˌ(���X�i�6xZ��VR�_n�C�[Ľ��*@���O��-
�g��dL������рpY����+$O�L��E{�t:y��� ��Ae�	ꭾU=����-����UV��M���O� ~۵D�fj#H4U���H%��
��c^�U�V@�cGc����/D��vXzL&�����W*\:l��(qA�a���e&��럕�]� Y��6�X
v��ķ�T ;��o���&+���:X`Q����v>�=X��;��� m�q�-��Z	y����F(ęF@8Ty��W*��:=�
�.hMJ}��}�ı���(��&�g�佄T&fF���{�,�Ĩ���2D%�rH�s�k¥�T��:��p�cƋ^�&�+��J�爡�BY��_���ѝ[�� �Nps����x��jD*�m�<$5��L�����n��`R݈bU�|U��I���.����3-7��Lv<O�y �&��Ӷ7y�"���!!RF���.�!`�Td�(�~��ɩ���kڅKa�	C�m.��!��MxPG[�����R ��*OVv�d��kJ�>V<����AS���ن�C�oߌ�	�X-�;y�	A6���ի�މ�ƪ��jq�͎:��k�j ��fa�NX�z��6��?}�I�Ϫ��f�������F�����c:���>6�g�_§�YԄCg�����kʌ'�ʏ��C:�!��� ��ȉJƥ�v,#��Z�A�f�aQhpF�IH����a��qt�2%��.�Z�1V}g����|v%w�N�Dg�C����X��,-�Y�bZ���;&]�Ջ��{t| ��U�տ��{��Pz����$?m,�BY�d�"=���N`M�YF�|�[���67!�x���$c^/f�Xtl?.%ૃ��⧀C&IP�������h��������('�]���Q�4߰6��;�,`l1�6��v30���<RJ�o|������`���>Tj]:�i~4�Æl��nM~�������)�ފ�g�yU	�R��4��C�.����B�uc�����>V�Г�_���
87!D ���v��Pҏ@W��M�Wb�!��2{�-Ye*[>��q&��cC�It
X�����e�x.�s��{�\<�k(�1m�����9VEZ��Fh��m��������~�"���s7��3�u�f=|���(�Ѕ�2v���N򾊍�D�ys���kVđ}��3��'�A�~	[}�/`����kL���7y��ԓ<td���n�"�(�X�f2�u��,=VIֱK���c����{��sV�@Xj�Ʒqw��'j^w�'�-Y'�ҔP/�k�F��p�[I�dΉ��LIO�FE���"{W娃b1l��R��J���V��ߞ�)O�����(��?�ℐЈ(���8�bV��p�`�a{���R��×���`�H��}��n@�! q����8$��n|S}4��?Z\���Ho�%�M�5��z��k�F,bk�<�(��9�ó�`47l?q�?l��6����%��|l=��-��t/[1��	O���-` ���w��j|�|3QT��&���K;�-�Пq��W.I5Lh?��Fx�=l:��l�+.~��;�0_�]ԭUJ#a�,:��Ny"vq_�~�6Smx����������;������P��_���"0�	�QH��������W7���� ]Y!ub��/)�8��Κ��0��B���PVj*'4u颂�;otE8#]΅Bd��J�PG(�#c�T�NU��'N�������8J�M�䜮r�9�d�\�tP�8*Y��;�6"�D�;�4��*+�l�L�L��[�4��������pjv��>]1��qS �m�5 Mjs�L��<v�����Ә���ݒի���mG[W�/C0};a:<�>(K�$�́��2�����:�����@�Sgkl��������*��t:4���J��ۍ̽��ú��V���D�1vۢ�
�˘Ė�5�XB���Je2��_][��)4^ѝ:������Ŋ�Ҵ�Q�
��k��3����ym�D�}����SF�H�Ur"�3�ٲ�'� ޜ6�+�{�t�
����W5�R�u�@ޢ�!���������=�%�d�6e�K[�';s ��;V�X?�v+�^t���/W���=fJ�����[j*fI?��Dß!�q�o�4�&e1�4I�~�鏰�ԁ����y'W�v�5[��ʇ��s+��m |
w'�%��\�����E6��F���x��w�����H�E#>�[a�E��꤇Keuv�	��dL�G�W��#�my�g�����W�k��S�j�w~?R�����o�%�� �ys=C�D&�GA/�:���x���6�6I���2���%�єG�oQ����ŏ�[8ms�7T��ݭ�oஂ���bْA@�N���{o[�1�����4�(��n���1p,L���S�~��HwW�p��!��2;��Q�ML�#���T^i�����n?Yq��+_�5R(g���0�V��(��XM�\�J��(�s?%����h(L�����)�^�Uv<���A���2U����E^<�~���4���a�R=|!���h%>);�a�k��E�tj_ڑ'�mh�U�����A�uA\v�y�����r+� �a�w�JG1 �`�&��0L�+f3�L���*�0�J�Fk���lu�eq����K+@hAՉ�s<z��?S2�"#9075[���"���
��^�߂W�+)���[�rJ�&��3���Cr�&�E�|����A�Í�3� Ψu��B�k3���\�s��h+�0ן��=0q��k����!o<
uR/MMY��7LO�P�ȭ��;��r���q��@��9z���n�^�,r��ܩsV���F�b.'1�޵�ڥޜ�;��vi�q*�^�xuR�H�>���ǽz��qu3�����e�����G�_}Xb%0���]�S?�o�Ђ��5�-f�Y��`� yørfx2p�e�L��i�T�OF��)�w���ʢ�j���%�9	��įľ�$��q���iՍ�5k"R@����\��\��z��Y����y�b�5��1�s3���\ qV�"���iѓO��*HwU��P�S\�@��Kx���%�kΕtq���y�#Қ�F��`�?�q�b�!�-�aLZ�;�e�AΛ*ˮ~w|��1\����n�<ov��rYf�#��Ҫ���!��=���������c�-I�?�߳p��)�s�M�
v�;%��R?ʸZ��f���$yC�ڽ]��}D�?H�/ ;N�C����Z,���6����S��[[G�F �Z��*������I.���
�
˼���O�7�J��b�k�c�$P2Ƥ�D��N��N�YZ�R8�mL�hh�������!`�yf?sv��h++ɽ".J������p��`Xe�-�k�e�i��e����$N3�1=8��i �ACIq��ث�?�|�F���
��>���ہ�4���5iw�O9�O���}-�?+E,��_�%��^�;��6���+�]�s��=��K2r��۽��w�¼�
����A����ӈ"%ټ������� 	˭Fv��� ��g�@	�ɏ-�_D�_�\�ܢ��TM5�t0a%7���e���J�ՄJ�x���4���m3*y�[e��a&��$����≯/�W��4T⌵���-���D�Ҁ���E�wfhW!��b]PO�|���B��bX	�š����a葉�[4Ԏi�'�������1\,��V��Yp,�^C[7�#�.���mMfP�$�/`��LB��D=�*�C��&�N�Μ�X�|]Ժ�����r�������_��-�B����뷊]e����켦9B�R �cQ��#Y���>�kB�i>����dv�q����v�������z�DA&���m&�+OW	�j�,c����9����p+��y�4�93o�ɭ��:�ra,Z�k��]���Vz��0�;&(��P|�O#j���.�������c�Y�U���#�^�+	�/C �'n����o�;iP̪��fK�SW}:=�b����A���W���>�%`l�N>m+����3�5���n q�XS&OȏDZ~�%�k�x�>�E R��b�(�ei�Okm�Z�O�,�Iÿ�q#�L�p{�rM��w��7ɯ뙽��ɝ�]C����q"������nm��I���}�� �����8^zr$�:��V�DD
< \��n�L[- �?��EW�ʸ�m�݀� ��&��IW	�V=�,�Bkl�9qT���웻(7sK$���]h����ܛ������+`K}�Ӑ}aOCmk=\x}��hC\=^qI6�
�~ӿDO=o����N�|�1��+7[�*�K\�h����5��/Q�E�0�P;�f&��n�%�g�@{fZ�	�_���'�m��L�[~�8ޜ7��#���^���k)���B^b�4�F-��gD>ĕ{�4��,DL�i�V.�>*Z<�u�H�1�t3P!����oi�������NIt:)yCƸFo����v�!J<S�#c�]b�j�.&h����ܷ>��o��F<�v��u�2є�Z͢J�]�#��Ky��#�t�!�Fh����)����Hk=
�'Y��"QȖ�F6w浂H/u5��
��ژ� I���񚑜'a�{m����B~�2<-c�!^�h)�1vF^<�kc�Z���هQ����:��&*3��X���ƺ��)�'��h�K�٧�1ivP�kx�b��u6;yK��=��)h�8�Q�e�*M,���L1�8�1�|sڋ����� ����1���ZS?�$"���A9��
����-hg3����M� 鯹0B�G.��ϭ^
[�Ƀvfu�O.���ӷ�����v���ϑ�(9� �o�{���I�H���H%8�		u���#�#�*0U�]]t	���ƚ͒L�':M�jn�K�������� Ҵfi�s��E�jDf0������a��"�gFϾ�B��v��IWϜ��?�q�\5S�3];�IP��45�m�|�J�Ou~-ݫ)Iش�-2,=7�����nq�4�%�l�0 ���g �u�݇����`=R�\(�˶�	P��bq�b�I�*V��pcj�����@�=���a�[	F����	�]��+�*�ν���6V/�J����c�
��V��ַOT��@G�������O �a�8�-�4$�e�eP!����kǫXJ{����o�i1)�[Z6�赅�W%ט�Ρ����G��yq�� ANQ6։D���e䧺�W�L\J�/v�Ş5�ݫIݭd��/��R��񯉛��m˚�k��`n�t]�5��@Lͣ�3����Z��^�t�*,n�w�S��������i%����*�|�� �&^�!�;��F��D0�i�z������Z�3t6�{�1佀J��ND-�aF|/˄!;!�ؠ�C;Y��,�\�!3#H��$' #un{�'ދ����h��-�6ǌO&�QV�N���8gh���_�"ZR�gR�&�|�n�8Ơ��X�����)����������'x�~�Ḑj�N����_�Æu8��pl���\����έ`�:z|���,9��(�x/�� bc^���Ӽ��F�8��ؒ)�<�=�k��Y|^ߎO�ظx`̓e8?j%ٗ���"�e?%�nϞpǆ����Ap<�IM����XL��ms�.�� 6�<%y�ɳzX>O��)�V�z>��.�Q"�~� |X��ξ�4�� ���"�&�X�����>ʣ+ՆB��6���ܓ��;�
h�~
��2ְ�����A��d�iv{ ����'�������O&�k��� ����r1��L��6��	�uh]�Ѵ*c�~��L���LAc�������p���yb_�X���(��i.��Xӏ��cN�����}S4�=a�4�Ě$V��L����=�L��� �	e�&��xGs%�|e(4��	[c\�՗��T�����f�Q�T�|'{@<9�6�E%�oV���Y����mZ��9%�i`�*�损�.��@>�n����Uz��T�z|�����{?^�I��1�j�i&�����#B���|�E�2�r��oհ�:8��p��8`�y=[ms|�_�5�������k�~̎�~p���c5���hR[��7��!F�BV��=sюN�m��e��)�O� �I�z�uȹ��,�c:������t/���l�N��[dy�v�v�~H|z��*M+��m�m�v�<��ٌk���$��?}�S��@Ɖ�\8d�=g'|)V�Cr�4���/�Y�)h�,���h椇^�2�kV�������N�m��͉����dc�_ Jo�����&��01hC~"i�&��ӭ�t���b���L�ʹ��ͯ�
S�z#f����h����@uut�)6��Mk�]a�e[l�Z�rc�!�a�{]=}1�gۈ詖][�(��Tc��p7A�]Z ��bJ�#Pn��e�}+�K�3�G�i�B?P���K �yQ����]��i�7^[Z\B�G!He��'�)u�L?� 6�B挿�μL_R�粬d4����kh���#���[�,��9��2���q��*c��A�
�̭U.+�����C����!M��s���\����b1��o(ȅD�d� e&x6�g�R����%6_z�7�gZ��8�t���IJ�<�z)�@����YFčFAF��i�2�t��p�{]ɀX��1n3����6�����쉔���&����|��8�(Ĕ(�?qզ�U�e����%-T��`��ğ@�nҢ��ǵy��<0�kڀ�ύ��q��$�{�aq�<��o��k��oy6� C�FQFeF����>��:��Kp�Mt:�<S����}j{�p"�ʾ	����=ThÃ��zp�a旮�	���xx�r}~�4c/��q��I�	O�# "�ȥ�L�)Ҥr�!�� c�Ȁ�=�B����X*��`���[2xѓ�^�I�u��&�HR��Nn��@zWVŵ=ns1�k�xCˡ,T�3�#f5R>Z��q�]Mf�����������ؔf͠��dH�j-��P��Hg&���a$��V�i���-2��x�d��t��(S4X�_�����Ú�Bܗ�x��z(�\p�S��+�n2U;�h8{�W���)�ɏw`�*�f�'����� /���hA��L��)5���OX�դ�d`�翛�	��\n���7%,侻�YJ}$��/�c�K�{�;xYc��2E���%������.m�a��~!7o�"��w� �avܞdh��e�e�2&��"�ܢU�,���ք�����l���0�1��5m�5v ��a�/�I�˄�m�f���1��3{�z!!hT<���xk�DKw?�q�m�j����ՠ��r�ש�8��F'_�����>!y���z�5,��Qΰ�vF1H0%,���XXƽV�ܷ�B�,-�,=��;Ĉ謉�!��k��i�� k����f�GQ���"�E��y�N���lɎ�)��ɚ䷹��6c��Yj��x}X6�~L�Y�e�4���*���*�[��4���Қ]���}�
���~ZK��0���7��4�w�ԏ��+�����/�nNk6�'#v[�P*Q��.͏���}�d��Nt���׽=���N[����	e�-T�ˏ�ET1� 9Y���q���Ȁ��ߋ�^v~�Dl/�1@��[3��h׃�,�}(ã���k4�����^���ڷT�zW�� '��j����-����1�<�S�9�`J�vC\ �s�{�������R�$�@TE�Iur�9�����`����Yj�<��fی��f�,vhd�S�&v9�Օ��aC3���u&�1�{˟<�DZ�v�A��?d�p�a?�׽dm�J�!�Z3%�d�/�+*�X6`d��U�擃W8DY���(��ǽV	M���n�A6��7g�o�X���YWMJ��&W��dK���e��d� Ÿ��G�.1���Np��O�N\gG��"�=�^�����x2Y`���(��pk���P#G�2��G�ԥ�p�v���rN2��-�Fd"��n��dW��t$蟾��N0� w"3�_*y���j�q� {����[�\�AcwE�?�1���[(����Z�bhץ����L6}wjov67H�CR���N;>P��"2�ln��Oʓ������B]����V�e� W�6E�oN�P�v[�"nY2fqņ�)��9ś��r�L���N�#$ca��fƙ�m"�a
���NJ��հ"i��F(7L�fª��_�0j�|�s�.��.B9JG��l2I�F ��h�˂�X�(,iv��o�H7\�A�������O��u�_N�I�]|��|tQ�WR���PUVc.�c�1Ǩ9��i6�BI��yݺ�E�2: YT16�3226�@�{�+���o�t�. �r.�>��y)�M�_WO����zs`�7�^��ī,�^� ��1�c� d�}L/�j�R��	�O*��\�^�M�ϗ܃}��d��˒�p�Y����w��B���,	��0*��G�{���U{� ^Yd��+A�Y��q��jlʹdTX�$[S����9���$Ān%d'TK�.%n��F����5M�wVv�P!J�a�PU�O�,��6V.���q�Av	:��j�O���{�b���~��d �V�ͽ�"[1,��C���&I�bi�\0�����1��6m��Y��HRM�ܬ枌	E`"ɤ���V�BX1��:��xF�����z��������	����dI-�{َ��J���6��j<& C�üO'�0<�����O0bzj�i�6m.{��k�>�I�E�������w�4�3���͏���*袑S
�,`�|Xw��L:Y>���p����&#Ewh))�����%+�ٖE��$��7DZ ��?ȇ����M{?@0�g��:B!���J�f��*�&#[n�Q���*lj���SѨ��"6x�.�Ѵ͜�p,L�p6n	���W����.�� ��KUU�G#�Z�$�|Q1�D�L�^��	����U���L��6��IT��>���s��{�[�Ta��t"�TWP�i��s&�k�!�A��F�B�\7�!�.���dGȥ�c@pL���>��Aڝ�E���'�i�"8�4���������� sSu�%i<�y�[ߣ���Fy70%�Q~٩������0�E��(��T��㉣C*OL��U���B4b'Fc͵{�Pd}!?]Q�f}ɻH��o��}���S(*<|jz�h?�u�3�L�'� ��`���h4|��լ
��LL5�����N^6�)	�610%��莁�� ��Y�%
"~M�uW�u�U¯�X���{�r˦|�x�2=,d��6���E�S9�9"^'O��4��� �RT�ig�
y�8IR�_�]�Ƚ���/#��P��H����1�K?�ǧ����fz�#3���;�xU��	<��g59VN'��ś�6���������&� r��v�λ�1?��T�6:Cb(4@}�ff%:P��<dIs�삹�(w�J%wtM4��e�=�����"�b?M�����N�X��*����g!���e4��}Q��N�zp��JD��>*�X{���X�߉ r���\��Al�4 \���w�q�#uyy�����knk�_��?���C�D����9�hR~1�z�?�t��I�T�jj���N��7�Wx�q���[��(�Z��HARX�9n���6�E�(6EZ�"���A!�T��]�g[�Е`R��G��x/�+��SB�0㹊��h?�CG֚/�.��bj��ZFOa��o�����
E�Ϫ��?�Ԃ#9��ם�U���n
0�R���s���A_�jȗh���\�����8�)�d�!eD|����\|�T.�!��Ү��܋���294[�-�CrBq
C�N������f���wR����~/��J�fF�b�Дk�*�5��L����!gx��9���C{���: ��p�f��q�Xa�Vx�EA�����"I�<L�'�q�C{�=����>Ѹ��sP=S�L���@1�����l�ȝx��Vs�L+�@1�x�j�py';�
$���r��zG�<�h�S���t�������C�K۞,J�1�Ȅ��,��莕-3dy��<��͞�Lom�<���ت�򚺱;	<�%�)ݐ��Ŭ`���'��<�ѬSc�+�mo�OY�����>�L�_IM�jA�Y�
tL���#��HU�~\/(nw=nY.9�9�d�ԥp�5����p!?���W��J&Q{Ŷ[@�ts��]c�9���9QO�I��XU r6�pl����8���F�~�3N2���qM�(u量H漲z��Rw�{���1x�C}X�s���#��ۻK�T�a���[Kd�����z&�)��!Ǎ|��*��7�h�ů`�s���Qx�v5��Z(zF���h�:QW19ɡ�G�OcH=��U[���H�y;S��F����=���,N���� ��_5�VY�7��By�r���;{��hߝY5�j���:�����	�D����J�fW�7��?>�7ї���ϐ5B�'���9�E���[?Z�Yzx��s%�6��1$�ؠ��G`��
ЭA��{5�P�%bu𵼺JS�1����q�9���+�UӗkF��,�}(�1�1E�I۠U�����Mf��)���:<�ǁ��@)��X �(���]���]�'�'K9a�g	Т�V@��J��~��i|��=�o�e����37�>��e/�G���>��z?��l��P����iQ�=���_%��`c)���P�9]��Vwȵv������d��%�J�!&"���=�C"�"<�q0�)�s�_��Un1��4�-<���kS<��5���KS-��X})��p�n����LB!o�F��YA��Mʺ ��̏ʩHƞ"�#
VTǚ���L'��X��<ԙ�k�zX��f6U��wѫ��;�o2� ��sy@�̈́.�HӠ�?�M�2fs��ح2L#_����U�1&ʬT�8K��sؖ�9~)��I�Ĥh�R�v���4��NO��'a��i���>��	�����4�SZ4�t�pR�ɂD�01���F����!'��7�ȫk}}��f�>��)�I�I�I'ԁZ-�5U=K�O�P�����B�̲
�5ctN^֔���d��֛D����pT�\�f��	d"�otu�fy�-���,��Xs��}f�N]:Q�!]����
�D5(��������A�J�B��>�w[Է	�Cm(oc�̤-֏� g/��̋�P���S�F�Z!)�rg�	9����8�Ԭ�� ����$�G?߈���`����a*xdGEҕQL%�����^�.��_���'�����=�:�YL�+&P��CY:>��ݼv)�� ژFSZ�!-���^+���'u� �!�ƲBв^��`���ƾ���J�����rJd�҆��I���hh��Rb��"�i>WC���-K�,U�]N��E]Nj��I1�-
�dr����G�>_~�2�W�ǳ'mtE7z+A�� �8��r�vWZ)�^�X(����Te���(4�Tޔ&(�P�xN<J\�|.�׊*����4�p�jE[t+@�L=��F��PTQKj���
/�<��o������dz��K����u�n�$P�p����F�֯
q�P�R��D�{l���!}�|\�s��ewi��C�ά�T��Zn ��7lj��1W4J*s4w�ŧ����-#߂(��_D�	,6,*��3פq}���-��@`hk�JA�s�r��	A��}l�4 M�o��],/�����4眥rv�h;	^�4�NO"�� vї�� �����a]o�����:m���?;�J�:��t׭U�S��W�� Au�����'�[�x&o��z^�~a�l���Wȷ%/QR;�F�?��
I�;f�m�:u.�6s�V�)���QQ�E�����N 3�/��ڣ. ���:g���O��U=�>G�J�{�����ԛ%���S�C{+ͳ���#�����H*D7F�������)lM�!v{_[Ѷ�&�3 ��"�$�R��u"$�%��;�J�J۹�; ;<t����!�x���7��@4`[�O�O���$*� KQ�=�7�`Y�ʞ"�?,ۏ]=��WA]F3�ڋ(ۚ���ʢ��/�	�2�����ս���s��,�-����
�~�P)��9(e"���ʯ��chԃ&f�z�-W�i�x��n9�~^ca�*1P2�MlR��7�H�Ž/g0 P��
9K�7#o�k�J���G�M��A��1��}�8{1�,�)��˖��4�j}V��Ac�!����}����nV�N^����X���
��}'�E�$ǐǧ����ZB7�X&���荍q���a��k���S�lJ<7�����%�\r�1�2��@�M%��[ZkF�Ī�F�!��U�SK㮒����P\2��[ĝ�r���ʽ��AC6�=�%m�f�}�dEE#�c<���hs�B�%,uE#�r��S�ß�����Pb�3މ.�ނT��֜�k1K��i��!�4�5M��"f֑�W�I�J�L�~i�����mѲ��8sE�'�x�EW=����U�~�BS�	hq������sV,�^P��9;6Q}	�]���a�0~����}�U�7^ѿߐ�������?-�vӻ�G�?�%H}0�-���&�U�C�\�v69Z�Y�y~���6�)���O���N^��b�{��c]G��7�@5u�v5r��h[��AQi��GMJ)k���P4�2XJߖ���:�L00�'<���H#C����RƠb*s�QFX��O:�O+T���N+�����k���ݎЈg<�+� ��`���!�n�h�6�9G<J��/��d%���ƞ��a-+�vxI�8Uc����ܨ�-z��5�������9�<��JƵ�Z~���ZC�!9AO}�F�\'.S�9�ع(��8Zjske�	TYc�1� ����w�1ǘ$$�q�!���Z�ІN
��4je:[7�����eg�5�R�d� �1��3��	���)�Dp�,��pg.2���lf�o�ܔ�d�� ��JHE�B�|���+��=P��_@�����|�`z���-�lh
w��,������bh�D�lꁏ`��6�� a���U�Vd/Z���Z��R �$_/鋟�F��*�Am=0�l
�^������+6k2�q��fp�y���HYI�&��1w �t�? ���*�F���㽑#s�D�"��:��X����@��`w8B��#���ٲ�|�ȣK�������6Ď[ݼ�1i�G|����;�\�fxo�'Ӣ������#�@#`�zD���˵B�d�҉��&�Z֫"��-`�j,]{�:�%�����Ϭ]2��s� �҈㣉H/GM)9aC!�O�"�8# �TгW�':/�/�t{��[�����"E K�4�Pe��N��[!�y��b��L��X�/F��=�\8�f^�P,�)��2}}7d�l��c+�1BE.v|ŭ���D��vp�4���=�-�AoKg,Ҿ�[e1�kNV#�)!�!�����fV�����������y�o��!L����{`�[�bX�1�"pW'��=����a_�4�� ����}?��ϡ�Φrrtgg}��XI���g����@�!�QB�����7�;�c��?M� �j�*��*E�(1��#�I�d�E�'b�س�;�i��p�{�"���<so�kC��x8	FQ���eFsiK@V �S�����u�lm)'/�z�����C�96Ư-�J�v;<��Ǖ���_��46�Y��J'��fM۬l�\Q��?��:���p��F�DԠ(�mu��B.|��T5��>x�|ϫI�����$_Ի�Y�*��Şwĥʠ2NbeI^Y��.8�7��kQ��Y��������Ѵ����G���9�x��Ȏ����8�|�i��v,�m,��C��?�@�Qq#��p���olڽ[��o6���(F_��1Y�ёNZy�U��p'��	W��f�,@�Ϣō����ց��Y-���C"v۝�k�R-(O�����P�x��ևY%J~�S�b{�/�NU�3��C���F)s"�h����v��p͝�,B��y�O����kN%��#
�� Z���F�OWP1f�Y��n�i7��CAk*���:���p9���T�[wZ#���h����� ��#; b�#(�ݾ��e�Oߐ�x��c?|L$C�(RI�n=d>jg�'/���vn�ڃo2n`{��=D�17�Pk\��h%�M�{ /�t�Xy���E ˉH��W�&sv�(��({}˗#���Ԕ�1�2��K9H)�ԛ�+r�Ş��22�|�7�qG�Ҡ�.A,Nz��4�F�6�5�������:��j�#�zgY����n�jdi��ejM.�i�7��7,D�����;�۰g8 �in�";r��K58!�vCƝ
o)J�ATG��}N+��h�n���V���1,�6'�5�������*����f�'�P�4�kU�ޞ��-݅�8�� +ówg[?Ν��(*��&{����7
���D��=�a0aX�C1^�΁�]��d�m���ɵ���7O�.�֚��j�_�.�4{0�����n�_V.��R�b�$6[%]v5��/��@��%e�`l�J�%�_G�?R�Yn��bT������� ����� ث��((�ϴT����#+j���?y������[��+�]����=��������#d(�T���br������CȦ�1g7:��j���Bc.@*$����� Oـ�+N~�B��KϬ�B��O�/��K�X�<{fZJ�0�����~ƳLq��1��=g#���݅=D�-�\��oӲ�
�}���P~|dF��ɩ�2�z��2��r���	L��Z�Qˍ:{�k@���yP��[|�Xv�\x]�0��Z�s�{�@u�;�E�X�H(L`t1�	�!T�-��Ӑ�>:���b5�6(2/���Ɖ}}��\G'IX5������m�-�|����4_�i���r�	+�-{�J��〉> ·Gz{l������. T52�C[�}5����|Ԓq؎��`9����/#���gcSDɌ�0 ��Y]�SI��ϊ��YJ�$X�咨��MJ�Ħ�o�D���X�!5|,��;�pP4gX�IH<�h&(b��I��1�������(<�®|bn���k��}Lxr���A�^j���wG��������e�u)����L�f�O��[�����&:�����pQ�'�ƈm;���RP�S���~L(���k�����j����Wb�!-�@ƾ��̈́�Z�`� T�I��쯲V�*��*9[�$�TK����2�5���c{p�VvjF$���^���LOԣ�)���*���-��|=���|�V&�3�{P����g�J�k�oѪ������M��<E|I����pM@���ԭ<hy����t_�IS��0,.j��)��t�"�|���^Y��n'�5���QJ���+G�u��Ct�����W�p�gu O~�bp��Gz��w��/P�x���͆�����8}�a��k"�%�ۀa�Io-	]ڕ��P3l86G�s�I~�"��/��.��z��ۥ�J���8		��aWA=A#,Ped~A49]F֖��,����1+9�N�,����hf\�WY6��vX22��Ц��h/J��dK��n����~�f��ʨ�7XL+O Cc������Igį��7��9�&N�U��kw��c��a<�˭*��~PAρ��O譠��#�m��T��VX�����F��[���a�
��̂�aB�k	�;ل�%ꏶ&����h�׊@�����K�.��R�7Ӥ�FwT���hǾ���
�9�iD�}jc� 9�N��&���4�����@��Cw&ז��o�6$x�n���]E>{�D$��0(�<��+hG�avCuP&^E��al���r���s��ٲA��U�.��wl�ؐo!>)��H��,��{:"t2���3`k,`���N�	+ }L�ƟǨ�AY���]>/���<@&�=t$�F
��_�b��O�Mx�e�(��X�H���f9�ڥ�ٳ�t�����p�ؕ��[R�r����������q�;��|Q��,%�NT=�z�ff�<!�Z�HM��7-�GU��~O_n��e�%�yРҟ�ed}����y��q���}�ջ��NVS����@)���_�y�{�!�ɱv� x�(,�Q�c��~s�ر��9� ]V;�G4�ҿ$�$>���]�u���~��`P��1I'�g,��)�v�Q������%��c�G��H���������h����8��aI��,:��-%�r�Z��㷕��@8�n��V]s�a����b!�����6@��K��^���(�!g؃�{�������l�Y(:�Ez|�Wi9wcCG�c/��|��
K�}������	�l[���L�J��Ț��xTb<���I���P�`�=3BxM�1d�Zp��������)[�.%a�A&���D�tg���?(�DL;�_a�Z��s�����@�&;qmI��t�����<S��|�����`i�p]��w����M�YЭ�2�>3����R��YU�b:X���,'"�G�ȶBU
��h�� �y-$�+���?�6����'	,`˻(����x]`(,����*�
a��;⒌�g��J)�\�r����n��n���20�C���
\���$B�<�?��W1�q2���b�с[���<8)f��_�9)jO�sۚ��Љ�hO���xQ�8�(�����,KC5t�y���0�
�J���������p':���5F�%��:܀�aDa�����,]�t8�&������٩�:<���a�����s��:���}���g	 `�+X�*��3at�gg�{�D^��5͐�^Xʰ��kEF�)%z|����CE�X-,��;rsN�sM
��5G�'X�9��FDc^�(���!�JT=��-u��C��'�X�ҮOaP�	T~�s�6t| Z��_b#@[%9  ��������k��
z��
s'�RX�dr��`��V�(,s^�w�r���P�H����?3�:a4T����kn�Ȗ恉7?l���Dia"#�Wp�]P�m�)zZ����zt�oH1�v���k�]���o;��RVN3���l�셙H��o�AgI��#��q��S��W`+�q�{1�%�OJ�Ǟ�1�У��~��l`����F �3]-�]�I�Ђ%�����)��n���́����3����7.�G�Bn27f<Ҽ2&��\sKj7������zh��ֹtn2�MU)9_|�h���@�$0�߆��sk�{w��N���
��&�iI}�B2c�G&��Ξ�{�BmX�i�e��J[vR����̆�c&�� �*�9�8~���r��x���ul��o^�ﶸ�!p�3�'� �u����:��Po9S���~�;D˒lN�}�-���%�,
��*�땈\8�[�Y�O���t�Xs�l��u"T����u�[����r�4i�A��vY�ˤ�|r��)f�j��6�|Z�� ʎ��7��O���us�l룣�n䝢K��Y�"��t��YJp
���sn�ސ��A�e+yl���7c�N��A�\ZC&�������BdVl�³̩��=�wQ7gJ��$�Ɲj&�Ou�H��³녩vrE��?]����j�ࠥCA��zP?j���9{Or��eڶ5� Z�&PZ�.Ư��.�Jᔤ<|Z���*�eTva���FpD��ml����<zʊ���ܱ���O�f}4���I2�Q�\��ݰ�=��C]я�����]����8��~�,N���C��8�F�G��9�{{�����E��Ô�Ek�OT^ �J����lw# p��(o~}���H']Cr':V�A�U?�<}(�
kKnf�C���u��.��Q�Z���k�M��e��+g��8�}��eCE�g����ؓv[W]{��|.�L$a2�gg۰���5�"D�<��Ee#��I.@��u�(=�;W4	[�����H'����S�g�ωP���ZJ�ax+���gr.:�]��7���T��}��ˈb��kұ�!+�[:k���[�P!;m\��UNH���бsY
;^2��Q�)���������\i��adV'����zR-����;QS[�2*�&�}��ReF�D(��gs"��8��C0����D��4h�W�(� �AD�D~;.%�|����~�._K8�����������IF��;w§���C�<u�y��y�&�Ѐ���Y����N������MN�"�R\��p<��a�3,
�薍u\�j$� �����Q@D�)�"m�)޿E�����������d���R�$ MMϥmF�{e6�U0���Oq�ɺ�8��;s#������w��l�s�+*MA�k���Y��?����DȻ�3dN�Y�m��0��&��?1L(\|��d�����ׯJҎ�xc�B���>z5tG�uuFE���]�/�����P�,�4p�7C��f�jk�Y�"}��<Y�]E�f@zƴі�|�	��㻀��-oS5-��A��pp���r4n|��l�j
��j
T��	1Ƌ�����-^3n��B���3�av�;UB\�|ӿ���y���hɎ6�/�m~��H}�"u8e��ӋK*؋�ia�!4�#Y��3�_{�C�9�!�1)����S�X.��۷-���f
|JK�8�b
�+�&[�%s��+�$�a46��,!�e�k��\�{��{�7���s�yHoX���/+�@^a��g�ܚ6h���Rt����*==�ub�|z,])�����"�b��X�{��D�)��" p��L���骧���@O�!p˸�h6 �8߁)�^O��|����)�X���U��*�6��?�9��W?�e0!�-NE2ؑ1e�iU�W�����y�ݧjE��?��>�1�yO��p�Nd}=G�M&܁ 1N%�|���j3�����n��lm�[_rg�
�D�9������p�OBte�����$J�j��m����XF/~�Q@�A�CB�.��%�����(༥��y�>Y�_$̛���E�o�>�����,�o��n�L�3��[�
/s���7R�n+.�{|Hn_���Dj}/g+��BN���J�r�rRS)c�G���|�qN�X> )��I�c
?y�#)���_����y���d8#I}P�:@b��Ku��T�zݼ� _4�)��WѠW
���9�ч�W��� ���xp�e4�^���-�;OIf��C3���6(5����CR����P�ֱ���q�[㌣���^)���T':�P�_���"���#8,�[�2��bZ�Srh�8t���lj��<�4'qC�Ԛ�O�O�U'����)�����Z2	���x{X�N,�P������ ��6A�#����V��AC��x/Q��@���p��ZI���}x
�ޛ��];jg���Fޝ� ë�W�t	ŉV�Qr%T/b4G�_|�'��Z�C� � 6����0�y`��Ə��.�O ��76KP�E����{�����s�D����'r�t�O���׸�?��'0�o�0kiQĈ�ts��ҡ���]��엊�@�T���1�ʨg�O�&�yԌ8y�QVZUL�����PZ�l��Հ���66W%iүl��}�#���	x���p�"����,��K�1�~�]��B�R��(�VX��.3�P%Z�/�U8�o9���6�
���!���&<����m����-K��s��s{5C �z�Y��8�/���G��_;�jT~� �0ݚ�RYV���RyG[�m[AL]Q�1�^�g��p�x��*tn��r;o��֨*�H�veZL����p����l�G���!m�Ns��'�(���d�6�=��]�Fn#���kLg�Zl��L(Ϯ|/$\�)��lB�?m�DA+��y�����\�mt�pgD+�t"�jT��
�͟^�1l��r�W�*��L��[q��ktD<p���4�T�~�"34��RJ�'8Q�d��qc�Z�O0�!SeV�~�iޅ^N��A�fk�#]���S�0	 ��6��=kI`�%6G��P3}|���W5�����.d�N'8V*7�o#�>֯o���jZZ�n �d4��Ή�UR���3����sY�Q�G'���L��D8
�X�{ڕ�?G%�*��L�(���	̾���P��9�s�Y�G���g���í)��:
�5M��M�H��v5��M����֌SkFg(���V%ć��h,W���>�3�\�j���>��݉Ŀ�4�82c��o�D��b~��£x�q�OM�g��'$V��x�*����øApЋ��F�N'̰�bߛ��<��ʳc�	2�;��@9w# �C�0眪ax����ݴ��z�-)6L�r088}O�M���v�g��4��2��}݌��e��Ԥه�w�b��&���v�#
��j+9�#7�v�j�Qń�T fr�f�my�w���8#o:��oD����m��qL�߭1=}Z���
��a]|c`�@#j��6Ixr�.Y�ܵ��������C#1)� �������}n��,�S$��{��y��V2���)W���A�I
����e��YL�hSGc^�<u���^Lⓘ۱M�����-Ƥ�����u�H��;k�����I��)�ĜX��,� �]����!�	�V�VGN�:+���3�R�Y�m���%������)�#�YyH0*���\��a=�Ʉյ0��F�`���Nf��k�(�P�]HOT�5���2tȴwz	�i�G������%ggN�Rmo� ��0|�7c��P	Z?>\����h��K�3Ww�o�(�л��F)��Le
��},��.������s�T$�o����3�l]��;�WI̿[�DJ�7㍍�ƻo��VPp�7ΨٖO���?��� �n;�GVkM�O����i��{����ؓ�]�Y-ں�I�1CDے~�TkH�x���Ӊ��GA[k�uj��8F�7���9	֘us�����>Idt�$�fǓ\u�`q'Zm��?#j��nl尞�>� ��F�ODcc���<��?���ƿ"��nF�	�VF=r�!k�D�4��ɣ�ݴq�߁^�OU��|gZz�k� ������z21�6�o_�z
����&���D���B�Y���N#w<z�XUN��0�Zu�Qg�FSfu,��땳q�/�x��H6���D>�5>�Q���iP��}xnv��Wb�[���ue5C'9�ۚ�2M�E�ˠ���l��W~ǹ 8v뵓��(�)�>n�D��D�s>Ft	S���{� V�{�5�6<@�Q�F�?�4��N*V��'v�J*9�b�p�.��OȌ�����$���S.[�rI[��ߕ��k&IҴ��� C=Yکڬ��r���6G�)��&٢��O��-3�a�[[�Qѣ}T���O�,|��rb*�m�c�F�=w^�(,d*.�(d���1'v3��8�I��VxQcSBp����pz˾��9g�PVȤ�m/E�޽�3��E	��\q}���=?��^TMsi��ju9�Ďֱ�X<��b>{�"��~~���'0u�C})&U��^E˻|���+�Ǩz���_������0�V..��Q��.&ϼ�V��Ï����S��j��^p͸ѐ�� �yt� �%�"e�T�� Z��� �7�y�̢��e�S�$d4����Ǯ}����|�7)�X��3�w����g��ܑy5ѳ��d-�;` �Gp1ܷL��H���T�ungy��n��o���^O���\<!X�Ş�.�Jp_�:{$��hL��Gb���PMfӭa<vC��n����JG��$-����i�7VA�������ĝःs9��#��H�[��W���"��@�xH�|õ`�:&�)��a�˝%D?__���r�n\���c��dcd ��{K�;�7?ۭ�Q��s�wb�)>3���d���د`����o�A��	s7���G�g}�Æh��I�R��?�dy�!�"�IE��+3A���}h��L��
+������A�H��c�����F� �t� "�d�ljͫ�	|Y��Y]�9��Ts�h��<KK����a���C�o J	�؝���"#@)���aR��۾%R�l�m�qYÀ��	�\�M�1�׌4�C� Z~m��aI^���|���b�g���\ߦ��)gɶ�/2~K���7�d6��J���5.=��R�e�6#�����Τ���y�OL`��h�p' Q��T㖨+e`Hq[�T�b��0������b��X&���������Z>�è�y+���_r�����%H� $�p�N[m�ly�^�#S��z��0���i�J[3a7��-P��6 oɩ��++ok��}MsK� ���0���_GO������}~6��eUT��]=3�Sf� O0��#���@ǂ�0����ȭ���gM�����}6I�\��0�����n�j4w�VK�ءU�����L�s�0���rI��G������"�.����`�ހfk���O��U�)>�L!+�T�Y����is�KE&Ǿ͛G��;{x�j�SsQ r��[,�ѹ�*Wg|?���� �"&�5�j���d�6�5|.�$LŒ| �kZJ��]qK�M���U��T������8eYՒ�K"��B�U�T��	�	х���Y���+Swq"T��T(׎��p�E�p\�cJ�j����w��l������"�z�D��ӕi��!�#N>�8FA^^\$�	􃴛�řū��f�lu׶��fbɔl�0K{�V����z�1�[$ze�@��R� ��Dt�2��lP�;��*�.�Y/��҉%��7�J�e�X�о���E�'��\��������|�9��(<�Ēb(�Nٵɾ����,Br��ªx�/�8NGǸ���$����ВT�(���q?��8�u�qD��ZK;��r��
�~c�RH�fH8�N甭�゛S���9���>�$yk�˖�sm���S�۬`~��v#K����Y��ēT;^���wyo�/�:��?(�ͪ������_yJ]Z ��*�mײ}��l̫8
	�3���"e����7��r���Ѝ>4������_����r���_��������>;<�6ؑ�eIKt|�/=��,�_�6�Ym�/��3s�1��#	��n{��;~*r:�i��5�֭��8�]3qo;c5�_�K���% N�h��@�A���M%rh���3*�<��:+�+vO(a��i�@j�ѧp�ڏ�r�<;u�r�sw��"�Aҵ@ޙ�Ib���Dx�m��U���=�vN	���gn�fH��Ԣ�lU��?T��+e�: &f��+��Fq��v�z�[(���T�A�5(���ql��t�/| �Wn��mF_�oUjť��q��$Y#4�N���i�,]�.����g*��]��ÐN���˻L�K�}�
�s�S�_�>]�!�@���G�����8�4%�q+#F��8yPw;�<��M!��hWKlJ@\�6�.h����q�����=��P��##p�O@�6ܚ�wYuG̈́�f� 9��/� a�L�k���^��\Uɺn��Z��i�q��үM���J"䣘@�ｅDmƴ�r������-�U�b�Ѡ�Y�������O�wZܧ��bCI}e��[s�!�D%��l	�[��gv�جT:0q8z�D\�]���:�W��"�[,�6D����0�)Y��d���-����O:7���x����q!���lH ����	�P�b�{B���TD����G��f�>���'��Z�;=�v}z��kS�-^r/��怡[��5�C&n/�����P�����C�R�x��\���e��[��UJ��..��rxe��=��M�5�S1�׉*�E�T6/V`���W�PcNnH�߲pLC,q��\�g�zsg��=��ʷ�+ �Xw�XYe��(!Kz��5�7�R"�=���,�[\� �8/1\C�U_m����/@�%B.m�����0k�)79��)�ӓ���pz0@��%}����ַ�A�^���
S�*��B?GŤf���m@X�$���5�em�B�i�&Uz�;=H�����6��F��sŠآ��s �@�1B�����<q�^p=�a�+�E������Y�Au;�H�^��"Tb�|5#���ѝCmЭ{�R�����E��x"M]?�q��orz�@����(0�z� ��S�K2)���XU�Q����o�kC:�D6��ӥy��XC�����N,�(�utg��UWht�M��1�$��G�vP���gT�_b@���z$�SVHc��9e]_�<�e�j�I�`ʬ����Й�򰯚�����!s��jA��J1P�`�Ҷ�b�����,F�&�O0ԐjdEGzDo����c�������0szyC�b�,A��i���hmΟ�Fnk�ڹ��+�ɽK }Nc�ℸ���bp�R�"93\ee)�GF�FO�ޥ���$9�#�B��<͙>�9zx�B�q:	/�K�1�vdQ:N������Ta�����;�L�����x�g�WAN5M�9���& �̔A��[����&��z� F�^\C����cFVL����ʡ���2:c�>������L�v���/ (�*'��:��UaęC,=�+��h��qe�{% ���!�Z� |X���uAqǵDc�"'>�A?�|u	_���½#����8#z��,��|�>)%HS����iD�"��1��#ɸIS
�nH�1��&�9��Ǐ4>5��,�v�6��+e2���qx.9ۧ����RQF��h����S}+{"M�� F�vi�$�����#�ņ�#�H2 ��n�KTr��p� Z���Q�uJ�Jin!��A��$�Ѧ�L�$m�M)b�G��PH� �I/���	zV�b>�ˌ�z^0�Ļd�R�n�bBT��<W��� 钨�I2-��*y��)Df���:�����W�G�y��T�
��'�[ōfl���0�*�M��_Iw�rj]:�J���ݥ�=��2��6"!@f�3(�8��Y\_���oՔi��7%ַ���%�[��w*a
��:� )�[��d�m��H6���ݽ���E�1�RC1�a��o2��I�����2��*�zÊY���D��k8�@��4m�	����I<%e���h_�>\4���=�=��	��%�i�̦~��j�'3�`�5�
W�{��1ā�չQ��PIj�NƧ�Z��ŗ����K<I�)a�`-���͗�S��W��RY�hMY�zȼ�x,�i>���~�s�pU���T||��o�bT�Q�ni����j�.���'4Qu{�Иf�Xͮ����&ҫ��g\��>y@Z�(��"��y���
���lS�2��� >7�1śyV��~�M�e��N�|��FۻH�����������驑�(�M���eH�oUW�U�lkgF ��ROƈ��ʠ�]����B��}���7&Ӽؒ��8�Gr��T��Ɏ���f�Aw��N���?��dc#_J�q�
{��gH6�	��4M_��Li�E}ٓ�=rի�I��}y�)���y�����쪵�b�����H���O�& �ܹ��s�$�d��ړLRL{n���(0�Se��7�@��y�[��-��(����s�MɆ�c�X��sS;5���*����8�*�{��/f��`3.,.	i������O�{�p~Ak��u`:;��^���:$���t�T�OXne�_���U�/Y�ν��^+Ck����Z&]ּ_�\ �J+�_��{WI#{Y��K����S0$���O�%��$8�3Z�"'�7���F�p,�� ��oRq���^��掴y�FL"tAQp!B��7�v��^x��<�q�-fM��[z~�oR0{����O��i�F�J�A*E���Gw�6t��A{����la��F"`��~������z�B��Ruq��]|�ǭ)�i{M5������
��=5C~��\�n6OUU���di/q�<Wd���o��#��ൂjL���9�tW?]
4��D���9D�`>����.�eQ:^�Y�EpiD��	��R��1��ic�c9S�n����{rFiw�*)�Z�S|��d����i:��:؁��}����*�24�����2)�?�t��o[�CȆ	B��Ұ\�����87#�F�N�ZϦ (��q�ж�GHE`�P]�?>�Ƭ����@n���h�<���u��Ȼ�Ø�pN�]!�"ʎ+~La���gA�Q����/�6f�k�v�����
�Q2���x�3��D~��($TGM��\�����o
�buٲ��a��M�n����i�6�$��Z"���fa�6��Tߐ�`��h��'磓��[�W�e�V�4�Fe����K�W'��A���$s���lٕVE���r� �s#aa���k/EK�E#�x�=��_�˴��p���N_���H|a�ck 5����'_�`��MϠ�/ �+�<z@yi���na�>�ӳ
��g�x-�T���=@�`kE����`��zh^��%섥O���C����!���e�5?��2�]�'������ڎ,��A?�4w��^j�[��{��o�y�J��5�%,Z��9���\U�w�I3 y-���ހ�e��2qs��b����i�j y��L�i�֛��o�%���z�6���ou��<8-�ĥ�/�	���[#~ e�?��������d�3��'-�`��
�[(�y�v��\���qDXY6Ğ^��K3e�9��=خ=��B�0c�^�׫�%��ӻq���T'����~ �5s��O:wd�N�Fm$tӛ��}��Sj�/{rz�{��7���ܬKIqTUZ�-l >R;v��~�!�c�`ы�x���Lo�/zD�;�{�~MI�g΂�=�1�BIi��f�?]/���.�#'R�@�"&,�厔d�J�ۦ����Q��e:�r��gV����Na�p۾�o��.[i=�IeDC-<�&!ឭ��ͣ��L�(z����LX�U�M(����.�5PUɭ5w=B��`��󻆡�{�x��A ���9�.�.2�u��M�h����N�o,O��`������Z�NW-Z�WcC���s9F�NK��O8f�f��8u�'�$�@Yu��,�/~��!�i�]j��+`^؎n�G��"�*�]�r�X����SPn�-$nY}���nS�U���[�� �5�`Q��Q�f�(PF��9�N�A78��7H��gf���`����������wͮD�bO��3�?*�Mɯa�6�;Q3��+R-��t�rj�?�M,�%V��VO10�̆��OB��1Ai:Ǿ����4)�q�s���T�ȧ�E�<ʺ�� ��lߘ�J�p�v`:zΨ1�t�.��<w����ɫś~��83���e)��E4Z��Չ�v[�Ǣ0�%jI!��C+�����| �~�deS��M�[� }���=9Y���Q?�R�Be�6_���8m�Nߪ�����4e,���oU�ظ�n�,��].��a�ж����������hab�Yv�!����-<��7�z+�����N��0S�o ��DS�g�sȞ��ii�[v��˴v��34ĉ�*��f�O�� \v��6VS1ݘ�m:��R�:���ִ݈�[8Bi�#����wh��Kr�c1���s�;�D\������(!@�_�"�z�8�,l58�x>��Q�z��fx"^K�1 wU����i5��df�k�� ��2�d�~�(c!��O�(F0=�4ޏ��T�g�
C<&�zJ zd���fe^<��Dñ���V�u2Q�������F� ]D�XGS��s��������,��R�&��7:��(��"e��g4��� �)O��\t�]�#V�R̐=�����r'}�"������T�[��ɍ,�Ug3�n�*������ �M;���cV�ロr?-��N��Z��E^�w����
W�����.�:/���<[������v��}�nn�&YX��v�
8��2Tc� �]�$�C�ϔ��b�{�jE�`J���	�u��0YcX}������7�6����u+�h�,�9 #;:G0`���
|8P�L�QՀ�_*�T�Ҕ4r�B�ֲN�=x����_�� !X�eE�tǇ�����렿٬CB�]\����,���S��ݠ�LQ���V�Ѥr������<6�lrY�0�TXDꠌoV�'�H�h�c�*\9�@�n���ݰ�%���u�џ����0�3뉠1
:����i�{uwB�Ks}�ҭ��=V�9��VZ#�>��G��-�<��صoyklڛ/�\�`����t��I�5ۦGu�m|���� 4S��4kQ]FU7\�４k,�OuB��'[�!����6;��I���}���H*)`�[�kh���y���*�T��ǉ[��au����A��](ݛ�O�Ӎ\~��N��18�GL	��Z.&���=ǒǍ��O�l�)G�3!p*�[�{�ʖ�JeU��>�4Uh閷�
h�V��:�h�b�*X�l��[�(2:�*��Bђ���$���*��+Z��UP�;te�nA���煝,��P�M3F
��f�=�`�V͡U�Ū�1x2 �ް��|�y^x��@�P5���Ϯr�����۲�>��[%��iXH(f.��]�fwK�ĉ�_q5��ɈXի�f�/�$�| U�����؟>���,��烥Η�^����X�#vI�KZ��2� �?��u�>SF�K�s=�9Ss���w�=�Y�)z�<Ud�1�Tn蘢 �-M�1UhE�Ts��OE���fuC2-	���/v0ѯ���G��-�G�+�����,[��?/D���>�*S����s���x��@�ݷ�����צe`(p�{��y�9��Z��wE_���P㹚d�=�"ڔ�X��dlFR���@mm/%]�v��tN�5;+<KpB�������I���4P��nq	����5*��.#�IG��.GK�=vȢ?`G��X����QY/�(��}�<��T�(Ԏzp|��U�3�Чt��\a|Gn�1�kS��#�����\���5���<�99	\�jW)��LNwP�s� {zP6�.���~�����;���K�)�ֲ��ˡL6�ʟ���HK�[ ���]��I�cS���"3�a���QD����d}�ߕ�Ω�;�Q-p�|f���(!;�1����{1�2�����"��8�}\��NhM��������s�N�'3wS�Jl �^�kο�c#.�l����+n�jD%BS]��Xj7�*�Nv�%n9���$��R1�Y/����q����A-����6�X�IՌ&�yOQ�bDB�2fH��7�dP�ks���.zE��e�!t��CRxv�"���9vO�@j�Ih���/h��������/�z�������]����ك/�|�Q#�6�^�4��2T�;�q�h���Z�� ��Y���`:}TII�Ⱦ~Lh�Κ��I5.��M��F.��U��tO�q�,�Q|�w"S�)��:���!��C9y���\
/��6���k4�7�D�Uڡ��o��n�oδ������в��\}���G��	Zkrn]
4�O�����ww�����qL�X���&�윓�4y/L�U@]��X���u�N�tY��gO5\�B����ʹOM�L�k��$.�䈚<�0����>=H���;��>ֻ���V�f`ؐ6�`�s�"��0Y�`�Z��Rh̋��E�zQ�0IMU���/e����W}%�Ŝ��O�0<�^��{\Hk��?Q���Pyg� �~��h�0�<��hy8&j�v���:���Ѳ�r����Ӵ�e{�%UeSZq��f�Y���TZ�+�1��i ca;˜1K��WY�
�k v�	�������3���r��.�9�zt��.�����l�_=Kޱ��*�^����'A�|����jK6�4�nLW�w�>9��FO�o��
�3�\�YEnw�G�)���V������q���!Ħ,J3k�����B۠����X�h6��Fn:���b�;�(�!�l�bn�����b��py5�7�������c�r@ui��{��NE��E��d̚I�r|<�Q��w�J?6U ��S>|<Ӂ)�*��l���
��A��Z�X�3���9�(̮t���ƣ;�'�[r	�}�����(���֣���'ד%+�
��Y�iJ��cr_�ȟ_o�� (+�O�Z:W�۾���:h�#t�/���kh���D�x��x��U�T\=%P��N���o�"�ҽ���or���nD��r 6����2�o~��ܯh�m��u	@&�ҍZ(�#��2��waW�D�#�b�:����
�vk͔\��o	;59Y_e���7�� RD�}����d_����>���ݗid�����㚿,h[�I�5EB�/�]b��=�A� '��c���7�4|�Y�����O�@�eC�2�K�s|��c�����.JT�$��(�I%/�R嘢�а����������7rcD�e�z�6�F�v�O^��l���M�i�ƌ��{�MH��f�R��RM!�H���PD,��>���d�"6䓙��b��2 ���]�����٧�DPlWt&����7��mUל7�@���s�ԧ�z]8`|���]�ȕ[R�� ��$>~�3�U�m!��!�֢�.K�y�;Z�o�����5�1l_���7}�2��2��D�u��>�,g�\��I$�R���.A�b C���PUp�]p��ӏ�W����C2����U�v��˞2LP}���&5�K�Y*�~qU����Ԙ =��b͂�֞ �CW�I�d6��-��@d����i����rPe
n�]R�h!!	�-�Nt+Y�u�I�E֊� ���+개���H`e��i�!��9�`م���;��!�v\{���j���!�()�o��{&�m�.>_yuit��E�Qp.y�%��r b���t�,�nnn�.���k�}��Od��t�ؖT� �O�O�j`o�OԚ�n:��. �8'3	�}9]<��q&�����y��g3����>+X�'!�Ш�< �K;�q��Ȋ�\"j~�ݏwӳ��!\���X�ۣ�*�/,�� 7p�#Ჱ�{?H}4!{f��xg��E�|��xQ`	Mv�n7�{�P,��f��R�6,�'�Y�g��Y���Ö�9��[��� ��.O����v4�㠟G7�r���cj��AR����=WΤ�k#��'��iE:��&�/���f7�������#I/o����+11��˾��])Ƥ�آ��H;h��ᓰ����=ҝߴS4���[56=߭ �����f������<�v G���;��p=�^Ֆ��p�@ߒY�V�7�����_�"���ig���t�fq�}��n!AL��Z�h��3/�o)S6V9���+�e�r..ݡnпYG*�3��ӈ��x ��'��Y^� �milFU��x�>ޟ���9�3��/:�y�����.6�B��#���tm���C饕$�(�e�����jF۰��>�.��|��	���R�2��d����4��[�Z��,�Z�A?��&X�$�B�m������U�!��<�ս�1@�(���X(�X��=I�VE"�a�]j���S�K>���	W~2��Ѷ+��E$X�M�[X�lӶ/���;��
K�C�D��B�?����f�ƪ#��)��Dǘ9�������	?���4�l�W���Rкd���Oa��&^)��8���B2�������Xz���
e�w�g�m�V���I����`ob<�c���u��sw�(b�d>fu+|���h���� 7_�^i�5�+��\t�dЧ笥��qW�tXN�W�]��A�U��r�����������Q�8�뢯��ik�?���
�C�	�DԐ������ß�s��<��:�lK@H�N��Ka���zLS�|-h]0����[G����a���ǼXWJ^XV��o���Y��w��S�K��M�v�;)��$���1���1uÔ��[��3��Vg�ŃW.�ψ���9˅�dJ�nczl� N�f�G�D�4FRg��,j�{5N����c.|�K�2\��U�[z�y�N�� bA��s�4�*���Ӎqiv�]�;��fk��
�`eƛcZ� (6�Lv&o4��36����,z;k~��D�@�ࡨ3��(�y�T�L{U�����=׾�9z�ʾ'�ꤳ�Y�3�1������(gz����BC���>
~[k,������o�Ԋ�Xe��>�%��@C��	�&�륄i�z����9H/j�'�z[9zi����6ʜ ǃ�~\�v:�����}�h���	�b0y��]a�0��oW�Om+56��"�U�!7Z��A,�}��NL��v���p��c[X�φ;l*(�bL���P���l�j҈<GKq�P��kg�G�����e5v�2زO���qB�k8��02v�m���12�֎4��F$�Qn��7�2���荽���^��E�|�|6�F�����r(�T#	����	�s�9��
�@�%�V�EϚ2�-���˩N������Mm{�����r����[�ZnP7�L�����ˑ�(|�%D��P��a����D'u�c�b/�C�J��Z�pU�rϒ�� *d�'"�w/v���E�����J�̼�4*؉��J���>����"]�մ#��z�^��T�j�1g錛c�~B�7 )���	Y���:�gg�o�޴���P���Yy��6���@��J��m�v���}����R8��*D%��h�������� pK�(����@�{����4jp1��H9�ͯu*���4����GD�b���P�kC����3,�Ã������^5�j
`�$8����A�Ek����L�-�
�.!7#Krk�4�Gd��g�G ��(��j�"A�),MH��{E;]��&��-�<+r�6�����kǀ�"�0����qb/�g��}�˪	x�Ֆ{�8��5�uC�G��6��=��S(艹�ۏ2�����e�Gq���h�s�d�46�W�I_7��ڋ�o�����θŀs/�w��IЉ�U�[��Sg��(�H�����ԽV�ݼ�GfW(=~��Zk�p�KY���1iH��o}��텨Q5]���w��H\�+ʪ�ٔR��>m�e�W��F�h�G����A�_���"EH��*�~ia�=E(���Q~�6� ��B�=ݰ�/(ϱ����(X�-�ve�z�{�EM(�=sE���O�����y3O?���i��.�@m�'�^�q���&�LԤ��C���NG�{�w�6C{z8+L�Us�*A%���>�\r���Z�N�����_o�Lg����hZ��YW�&CM����F�]N�������O_�on��^c��;�T:#��fT�T���|/�<��/��cv�B��1�Whj�������cR�!���+[E��o���ÌZqZ�v�y��I��c|�����HhS�M�U���E��.\�(�����D[9�|Ѵl3���^���HƼ����m	!�b�U���V�	���ͨ�:H~?"!��N�\R�Ӵ V"m��)p��N\^�3{�4��)�򕝴�p�u�z��Ls}E>b�o@��Y ��X6��Yw����Ӱ�,�C��K�-j�盤��j@z�&�� W�9Z{2w��p�A퐪e�#�,���1۠�h:���8�O<@�_�yCs��g��h�7�N��Yϸ���R*��_(W-ژ�=�Ge���_�~����s\��+��9;^��xh���@v�٢��\��3��3�Z�D����d�O���QY�I\�Q}�;�hȕF5S�e]�a��D]qOc�s�`G��|�X-����g�W�ݕ\۪*�J�}����}vQ��"c�$I��p��V�(���Of=@<Ά��$I�-Q����w�xf�M�Ë�r�`�1�Lc�qH��������kN?�k��~v���69L����*UvQm�`�sg��)~4:��^�m��w���_)�v���w��:#�mͣ����e����|H�n>�������s?�N���j�𼃒�B�d�1}*�zpР
b0�Zi��Շ�Rk2��n��iVF��mm\(��bQ�����?����������%�7�k�ս�������X���Eh&@=@�w%]����<�=0J��E���P<鹡��}��ы/������ P�RO��?�2�ݜ9?��=�E�w沖	��.���j� �w���E���!��ɱ��8G�l�{��q�����`�uU�d�у��"���ʫ�h5�����B�Y�5��6�Z�)%��0�Q�N^�FD|���v�t��[+u4<�_����R�� Dj� /2U��8�3>0���_�{Aￅ�9���1�����n.���Κ�O�//Wd4���Tfl4��j�򯲙O�x�&i�:��Jx��gm���i��ku!��,3\SiX@^<8C���S\�#�G�Ԯ늇�q��V5�;�b[Tc��ν�Q<�L�;̐_���C�|� %xs��p��u��P�6���ܘ��'���s]㩅 g�*h�z &�%��6}_}!���;n��yR�o�W2_�K�9�p/��������4~m��p_�f�B���ൾ�c�K�U��?9񰈚>��y*�>p�0�����0vC��Ԗ1�D��'mˊ�*̕Þ�bJ��v"b��W�}����`e���������I��ե(1&�P��\�F�D�̃������,��W���r�Y
|Ɗ,=T�ht�S�9����P�Y��pCi)R�_�5E�!J���<��2�3c�#��:fAナ@�^����9>�	l֝m���;,!�_8���\p�Q6w��x��À�R��EXl�Efe??4���$��x���)�' >�a�+�tem��$�%�x��C��?�������=*�Q�k� �n5�*15|,=5�C��if�`G�6>���k^�W���uw\7�7c|�1Jc��<#�k?��L�T�B��_��v�� �1��·��M2A���?�@ٽ�)�v�{�!�����o=Φv�S�M�):� �Q?��h�XL�g���tvT1�c��s?~��l����D0ZU=�	�Ѷ`�ݡ�4s�o��n�Vh!�iZrR�}F�9df�]��)L�2��+�*zb�g��MF�K�����kag"�I�4�](�b�/&�J|guf��J�n�y蹈�Gٹ� �I�˿�C�����}�Vbl_��qO��c�g=�X���#-CLw��}ZNr�l�6��2Ci�# ���?��N��^3������EL�jZ%V	&�d7A��'x}�ȿy�3bTٻ�=�l<�xwDr0lZ4��a����ښ�^�pN�2M"���6o7�tɓ�z�$�����5�l^Z;'��K��`p6�s���Q�����3�)ݠ���mH�2�Ʉ���[Z��=��23o@Q�G�'��´}�C��]Jĕ8��_92�Ė��F�̨=І�OS��_�9�v��4��+��Po�It�4z̧���gҼ�LӲ岶:�d#�� ���ؒ������@ �qN�:Z�"�ux)���Z���LXQM���T��[�z�G�~��k��7W�����F������F�OwHuڧ�;�>tя��,�%S1�����v����e<�0ά���u�uOy;�k�'�C��C�t*k�7��#�b�ۗ.,�@ToG�-q��Z�ָ&$"m5Jp�-k����ٯ��K��h��\�Է^)�������i�(ZV{�}�zM�Riϊ�^�H�6[x�� q�>�^ ��Kw��S��fQv�u,��8�y������Y�Y@=��ыs�����
��������bG��L'�~ԻMK�Pq�^��k<�<(�	 v��de�8��eg��	��5���OL��V�y���,�x���NW��8��)8?>�R���D��U�~&<ݼ�zm	a*L��j�z�pg8
��,�5�j�` ��7�O-�=�����a��D��0���58��T'ЬT@��,B>��V�^���\x�����1�=;�n����e $=s���$�g�ab?��c���.���T?2���=�=E���H�^�0l�_���V-~����,�κ��mQOYĿVy^�U��b�B�緷�?X��aRAuy�D��DX�k���JE �����VW�\�9`uM̒���eÐܨX%�O������Hq+&�(&�s�^k�S�q��i�V�+�������8$� w�����Y�w�'t�����Ds6���G8��V<��p��7��'�U�z|=i<�g���H&ė���2�*!oM�m*�\��b\0�@Ȃl��i��4�x�M��7'$J|�C0�E땘���B�B�|n�2�S�����3U����}�B���(�{��M������[��j��Q�^ܜ#Č\�m릜v1����3�.����q�8F�n#�S��O|T� �W2|��)Y]Ֆ�`9�%�V�@Dх[�~����ҳ���"�L&�g+."=s�nϖp���i ��⻦�+���s$3��~0������Eٍ��)-((���CÉN��N�,��Hޭ�l�5M�i���&<����G��3�fm��j�<-�r�"#z�`���η���;��J��EΝZ,bw)_S,2���O(1�Θ�\�w��ڑ5�@�kސ����+�M�F��U�V��&P.餜t"��(�'�H�3��,A��Կ�+�%h���5�%���F��NOdK���}�g>����a��(����\��d;�i=����GCb�{$�����ݶq�lK�ܫ�.+�� ���|�����G��ޒ��t�h�?g{�"s���v���a$�T@?	� ߎP�WW�#�b��+?ҿXZK �;�լ�Z"����tsC�S�&u���#')y��&��rs��rr����
� �����BIh��n���)����z_*5c�� �{�&��	�F(Bö�`�b�xMu���Xc��`�n �{]D��I�-Ҽ�1O�s��H�����Ì���gq�$M%Ɓ��Dl�&���HB�2x����q�� }u#�u��u:ȁ�t���-Nu�D��d�@�#�&F� �+@�ԿBsF��q���>���{)�0���	���Pȸ^��5k<'z��~��0�H�@>ʾr9�D�y&�;[�ߗ�����X��"1j�GJ���Ӳ�Cg�w����8���Z$Q(�ZI��1.:ø~�dv����ˌ �pHj���EO#�o�i!���I�	AOy(B͈<+
8j�U�,7�=�l���8ČnȪw�i�ߊ ��d`)p.����P~�g�Z$VmY�z�XK�(����j]�!��r��B�0�L��]$�˙,7�����c�O�O�36�����Ym�,�Ѱ�����l��Ml`� �R���d�?�-X'�o6�u��lZ���x���%�&b�8�9+"\ilʰ7��������0{s�DE��&�%�e7�%~ $ڐ%�1����(�Kݧ�Ș�mz�v4#�5*p�B���ټ�=��XBf`8���U��@ຳ3K�
XN�=\������g�Oք^�w�r+�$�C+�&�o�
W�Z^��ET��,1������]O�Z��=V9-��!��(�X}�|�z�v���I!�7`��y�c�S�����a���għ�����x=�3ژpa(���3�=S�)q��d	*-���T��5�iyt�!�uŦ���Zm{�7 �j��c��*juV|�/j���nYP����+P+EwRI^ �>U���z{����89^���U��U�D�#�T)M� ��-�$a�:��G,���������R�`��>�/ɠ�т��l{$��NJ�P�8?�tP�KйvG���G`����쳼%��ԛ}�0��g�`3؁@�2:)^��L��������j��?L7�&	�b�'  �j?�7�u�je�&�U0 �D��^v�~��Hl���?����w��[!�.����jX�[���DaK��ѕ.#g�
َ���믇Au{^���``/)I�vP����aGZ���}��ǡ����yV�&�*Z��@淨_��_�h��ޖ�z�Nڡv$����%Nmef����ڠ~ׄݙ����ѽ�_2�7�5e6�gC@���,��B���-����U"�{��Iɧd�d5�9���ˎ�lN�"@�&�o߱��!"'�r����,S��_b�!z���{��$+&+;F���&a���@��񺴔�ߐ����w�~��J�u]W|��	t��l�\���)��$@�k,����8���S����9�.���D��{�u��H���J+�������-�oI�:S��o�YmC\:����z�yS�O�}؈r^��Pz�,9�9KT����""jo���%h�~ѳ�����}�	VJ�TJ��>ԥ-i�? j�ȑg�S�Oa5����W���C4�og��0�Le���X�~ZU�0������2�����R��s�5[ 
"#f6�c�ל�5���65	����"�
�F;dy،EE�/�S���~CQNH����꘠��Ы��k��z� ߖ�T��_�X�����$l`X��VMa��VekXs}޶�b���2�B=pM������0'����/g$d����`p��x7��j���?Q��Q��Z��y	/�Va���������ثҺ���[�c���[��.��2����,�  �{4�>��}Y�h�"_2Y�8��9�o�)�$Ǳ���0�YV$�<���Zc*)�0�@i¢�~#��?UWfcR_ˏ~���j��!�SI����oc��C[
�\�q�K�����8P��U<h�<�yֿS�����i�v���V7iY��5 =O��G���] �-jD�f�{j�2Q�n^�Ug]o�_��6zaWx.��#1�
nZ	m Eg��Ƙ{%�2jV�=�����6IQ=�h�+V��䵀C�65vY|�>}�J�_�4�����*qfϣ��2[#M"�h��	��Y�l�kE핮�Ý� @+���3�~!��>;�G� ����*�jP	�]It+0	))����L'�@v���U$C,6��V�HVHj3���d\kf_����^ff# ���"I��qpG�0�[)��<x�����DWN5#�-y�·_�\A�j�j�0��I �XF{quB��4�$���8��J�aH�RvJ��Eє-��xs�]OH���t?5yk=��RTWRA\Z �I���$h�R����i�4߸c\�Y��u,��0m�;�퍘�5"0��jQ,�U-I�S?�|�͙����ɽ%O�%]uK�P����
�q����H߆K��[�M�޽ J�s�Ű�VBQ�г�~�e V�mL�k"�?O ��]�[n�f��A��C55)�w�����o��B��s��p��i�7'�t�m=�:K�E]��w.���X���0�Fq�a�TyH�7��,���_��,x��V�n�Yʈ��S��x&��ǚL0y��6y�O�����`�4g��ʕo���SX��$_�̚%���f��AzCѮ�yd�����U �!XO�'�Ze�T'�0iU(�w����[F���]�K��"^,���v��u��Ȕ����bZR}Gy2*%�.�����'.x�.ң� �B��t�%�s�)��:�
ŭ
v�� �ۍA;FK�#�����.�@8�'���CR�_H�{I5S��-jΞixZ���I���`�3�X�5ר-�[������tE0X;U=��P����e�R9�Z��Vݬ%��T��]�IK�&�RYG&�^S�c,�3��za���j)?"��Z#�i�!���)n6�y!���oϖ7��+����ţp��d���5\��~�
�G@clߑ��~e�YDh%A`��L?0@�Z݇_7���v�u�Qt���d~��� ���~=�Q��וֹ%#�3�3���ʷ�LV"]n+��ʁ,�	��ݛ� 
6��䋶;le���7p�W'����9h��àn�bu��?�m�9�pc<�r����Vc,$��?"�Q/�
C�U�*H��S�4�Ӽ�����d�Ơq�����\���K�bK���~�v0��<ᖓ"��6��:�Z��+��>n<kg�$�Wǣ���*�S��ĺX��|����!�W EÀ��s�c ���p0X�d�?�BA<��O�I�S��-�_�N�5�F&�M�
�*���n��y�Y�Y�"5L�1�#F��c���M����p��1��:E��>��'��^8S�j�w�"�P�9!{�G�
�E1%9	�Q��PqmG��~�����$Z�y�첒��U��A����^�QәH�blhxw�4�z��T�֠cO���
^�`���8N�I6sˆ�pL�/��s�µ�B���S��-Oa�JNT�]�mc��k�I�ʁ��/����>��r7��ߙ|+���>|<=�<E��p��Ⱦ�$��A>ؖ;ʏ�}�mdaD�g�b¨�(�������B4���ҔQ
#.�`:�Շ}���������d��pw�Q�4Қ��_�PЦ~G�_��8���ĝ�5���W8�ǟ����C��ь�l�ԡݸY�b�Ȟ��$�y[2��&�m�w3���#�p�[.��NX���E3����n"P�{�W��0�q;�v�g��LJx%�lZ���;�j��=�9U�Ҥ\G��z���ׅ�:��T�`5۰�W��8XĹ�-e�LQ�#�ݜ.s$G�g�O��M",�s�,Zh��f;K~��a�c�?%�)���ԾR��v �{ �a�p����7��V���N���*�s�x%~���k��}Ew2`%���x�u��� },���͘H|A~��ۺ��RG�����h2�?���� ��9�߀3?�i��B���>��U�#�V�2AWW0E��$vA�bZ
F�V�-�k<U���֙�I�N�T���<F�9��}G��~��͵�>f��9d�pt�qqվ\���R��U��9  ��U� �|����gvg�yy1P4笂ى���9_T�Lk�:��u�_�r�W}�di2cvZ��m��_���ؽ�8��<�wR5�ob��S�b2_l+^Q�\1�7��X�[
��ҏcw�2N�}ϑ�ş�j�׏�x�"k�~�C��,7V:���2�L���F�=3���kI�� �e4�D3K ���8�U�l=r�,-!��޳���&,�_�a�y����*�_��e�-�}����@*�-���	~ʤ�K3 B��8Ϸ,L�i�'�J{:ץ����K/)�^.��]�l�gRQ��J�n;� l\
EU�1�h�Cb
�Z�Luiy||�e��$�a�KP�2�3'VnҳWV�L���[[^+.��rG���S�}��/�Y�:�#M�C-q��	f/>'����PLX�%��0@n3�b�
<F�L������7<Er~^'w��m��cn0��~[�?�d��3����*�8��=��7��EQ@k��%��L1���0:���D�b�@�:�M;E�l�z	vva�����{�%ب�	n�BW`��,�C��j�������2#�����`z`hG���S��u��rw�aղ���� n��7�F��V\M�S�<��@)���a�����C�Y�ɰ-.ox&=�ŭ�X�M|#n�`|_Q|w��z9f��f+͛r���%/��쭘јm��n�@���Gp��G,�b�q�Eାt���3ۙz.��%���,&V�x/�V�1�Ϯ�&�@R#�+��b�Ӻ6��F��b�:�6���O�ջe�?���PJB�S�sƟ�R{��w����`4����0ޓ��j)�MLS�^R䮬	�=mX�Z���b�)���!�h�3Р�)�p4��'�F]���-7Z��Cfа�~�H��|�ҼJ�� ����������f�BPj�!c��dM�8�j,?Ͱ��U��y.I�:}?�=c��k��)[�U��ZN��-���Ve?V�"�yk��Ϯ��Hd"T�QUl:	�4:��Za+{�3"3�O�~��A*���-q����sx�>�đ�x>	3��膆�9�)���s�cf�	뵳��'�!��+�B��#M���߈�°=Ϣ�#�0O�	w.��E�L���>u�V`b?f�)�P���0�F�&dB�����ђ�n�Ŷ$�c�o�I��0�����t���~ddf������>D���qӜ{��A�� 7>�\ǝ�h&�����JYs���z��·#yӅ�p�U����*Ϙ���*@��n��*6�Օ��Gڂ=AI;e"t�]�2z�`I����CZ�s���ѕ3�֓�{�����k쁙��O���O���.�Q�7%�e*G��t�/(Y9�N��3�>R���Z��ܧ�6�K��T�b�[C��C���SH����-�JǏ؀�۾�O�uӑa��f�}г�oU4i� �����M#��(�W�X� �=��|�]}d������(�`�X�Ƭ��%�y�1CN�Kz{�#�� )o�gE(ن�х�9�� DH$X�T����{��ߎ��p0JP$dْ�w��*PK�I6���'*ENQ$�4S�!��l:"�U�C]ƒQ,���HС;f-8�/�j~��j=k��B3���YC�kP+�#u���w�@V�]�j��X�U���-P�ΐoW\��8Z�J?�3���~���g	Dk�@NYЧdBw�d��¤�nQB����j�ͽ�I���R��*uP��3����'=�|d9R3��4;�<�?�˧9\�V;�Na�늉�/X�x��\<_�j�0bx�T��Tk��p�2}�!H2Pg;��L�@�L����S|,A�*JV��L/�>��k-��W�l�s��sʐE�+$���t/�ᬂ�󭇴7����AǞ����O���:�|Y
f�r$����]4�mc?[��Z�M�:��\�c݃�n��8�sӮ�Z���Hȝ�=>�d�hw�5�+���G<h�g5e�k/����� ��+?��{Z-*!��A���N|}>�kpq������8z����,�.�)
ǒ���p��}�U��@i-p/.3�C����]E��
�U6�����ن�_�8Y�:�];�М�����g1s �����m�a��敵�ϡa+�E��X�R��;�:ط�6;q�YA�rc\�/�/�_(�n�8�g����i��ݭ�nr�0�3�D��$%&K�N����	'н�QU��]�T=����|\4�kO�D�Z;$�;s�®��P��v؋�7B|��7����*"1�$;Vs�u%=��}��o�˖Ӹ��B9��^��f����_Si��9�}�.�
���!mQbbs��^:�W�H�l�L�j�6D��ȌP�w!�Q�={8k�	=�;.|�؉*��G�n 1��F2��D���`~�ʎ��/+���&�0��V��(`^��=����6vnۅa�{K{���C�<�cܧ�D���lv*݁�S�E�1b��hrF��_ik����U���f����]]ʷ�W5LPl��Y��K׼3�����L���t���F��e� ;Z��V�Dz��+[C�sV:eD�Ks�v���&�\z����E%#���z�4�K�"N�Ha�\b�邖Gb"�5s�����ߤ�-��c�/P�� �� ?7�!IA�)Z&8�lH�hz)y�w�M�%E��w��[d��޺ 8������K�_7�)�������:-PЛh��&��P�d29E_z��1����х���G��}<�a�񴔋��\��$�9�� 6'2"x���\�W�n��2u�����_BwF���գ���I3�#�G;�$YCj�[�D��
	0>n���⏵������4y�q��^6�L���5��_1g1���:P�D!�坸B�!��!U�	{�Ԑ�2�O�p@�U�Y�r����
��
��j�0lR��Ҍ�����J���}NIy���K:`wvkSy梁��K�Ŵ�C�M�z�Ӗ�H��;�,7��NE1������j��03s�BH���}��q����Q��VЫ��� LX4/��>�9��3a@V��� 
4u&���*�pXpD�n4��̭*��+{�|��[c~�hf�L� "6��Z�]k��q�@���is�{}Q���u1�k�0дtN���p�&3��:�T�?���C6�i���,��𢽤W�25-4�k��l��!�׾QA>$����;���.ˢ}%�J��E:���R�!B�蜷 W�?��S�@7���a��2.9
l2>���=y|���n��Y�2e������1T�G|nz��^ʗd4[>a�H.�(SP�^��֙��r������-�w�	�)3���/ew�h��S�:�a=��A��3��f�u�e��x�|
�i����!̓�Z ��=�o�v'0����w�<!O��ˁ�ngt
i|�/f�V�7W/Z�LMk�rb�� �z�L��������?)=Rz�3�@*��m�o0iƷ1�	~rI^��2�F�%Ս,P�*^�L|W1}pkT��~;���6��
��̶�l�Pe�I!����텲[ι�oCP�y����PU��Gb��>*�B�|��5���cx��j�%�?Vٯ)=3\o�����̈F��G�^r���IY$�XK5S_��c��S�7]X�y�g��n`Ե��Җ�*��}�i[����p�d�3PcMi׀\�Ǥ:|��p��%Q��,�[I2�Bd���)=lgM���MHE�4�ktEAO��27�Ϧh,�����?f�ҵ���0��:��ů�.�KN@�*n����R��*M��S�`L;�k#<9�5%	��kR�_���VXˮηWv��<��7���H�Т�_���N \d�ˑ���F)=%��`͕��Y����b��1��5�=�?�j��
����U��شH1��|@��GѕK�/�mW����ۄ+B��|�rRP�4���z@���ݠ6��0l[���e����;+�tZw����n�x֕+��Lg�����ߟPz�3'k�}?sW���]�5��^M'�3b���I�9"N��2XT��h��@��j��=$�q8�
�җb����$W����g�}�y�q�#��y�<�^�K��%
��@���y����0��z��z��ݝ��k̖�9���Z�����_�g��z1֪~��i��0�5��
>͡0Y6� �[���S��q1q�-�y~>�@m��÷�g�&���|3To����fT�̮���M���T�$U*�%�"��δ���=�k(��s��=�O�z�P� GqY��CG^��ɋ:r�Q���C['�a������qS2��D싼���y�-��uVu_�Og:�i��<�둗��J���{uYdx}-���Jc�3Ӎn����G+� >�0���-u��:��u�y�)�Ѣ�,c�q�q>�<`��Jڟ�E����چ�U�W��t����T�>�d�������&WxË�0�2�\�|������V!�h��T��ugb�S[ƺ������9uF�8���E�ZA�7=��A:v�@�`#����F�'0�A(�5�����n m:P���We4�|��1;
�%e{�=\]����(���2o4���.����X}�43/n�PT�u�w4 ��LS���kP���V¦�*���'G��-�_@���i=�Z�/����V���Ρw! �����3���YJ�Dq��E?|Me�hg�i�yT��MT��OߞtT75����Λ��t�.��$�Ê:|�TN���c�w5��eE�Bb���竅�.,jOaP{e�[Fʓ�?�:Kp�� �,���tG"�|��� r4:L��2��?t��x]�1�"�8��<�K����R�d�XaKٯ%#6�``�{�G7-BV4�a���L:�-���ѳ�be�/���=Q^r���+ S{�3Ԭc�ZC�ZU�����W�^�UY�43���D�	7��i]��p������,祩)ϼ-��R8�^v�֠(�AI^6���Âg	W�|������W 酟�`� ��Jm(���*y�����b�!_�C��Q�uDƐE�{����Ǹ����%�M&�@@RI�4՗�Tb�3��r�[{��ԣTzO�4o�YQ� �7��uݎ)�1�Y�#°��J��&�vN}�-j|L\�Fa�����Q��.u��Y�6����т��#
(��{�񾽜�+��kTh��Lk%�>���L��9Y]t�eA�w^�=��o�t�&�V���?:U L��#��}e��@���h`Z���X�Ր��B,�L����V=�zʯn�ȨInAZ�]���&�P�� C{Z'Z� W�)��,��Y�T�~��m,�j�6����o�l��$vA�#]6s����t�����x�F�k��\E��g�R�ؒ��w��N�	����$�݂��e�U�N/��Ӥ�e��ڥ��$HZ)�h���@|�n/�$d�w1~q�v9**p����E�m��p{��<	�Cd0+ r���O�&2�huh�\)�G]�Ӈ� ��:,�Ė#Y2x�PK^^7��$TP4�݉R_L�KyQ\��
�/��s��{*ͼ�B-�0:���[T�s��wP��)�����c����^���u^v>.�c�(�L�������҂�i�C��ϐpI��n@�-�J���27�/6u9����:�vJ��g�O}��jP���/�:���������e����N��R�97��r=���{ݩ~����ʯb9�[����$�h��Ѝ����V��BϿ���JKh��5o+����ZY\ p���A"�����t�������As;�2/7����1�S;/�����L���&��$a$4�ė9k�U=��l �JB���.��� KN����<+�'����##��&<�}�����ɫcm��PJ��0<��^�.���/�|	cY��z��i��U����(���/�S��F��ɳ�GqS�k�*�.\%���s�(C�#���,� ��=�m��e�w9��W`D�AY%(���d�!�˵Dׁn��U�s����;*#A����Iu�j�(Rn����e��i�~v��#Ix]+bIV��9�H��Z?�/3��/m�?4�$N���s�J��~
yé`�ہ�v%��y�q��Ҥ~x��o�59<��(8yIO�\�}_g��`�<m�F&��he���%\ĉ\#��_�'[�������|�Q�|��B�y�V�4�4����'f�)!@�Z_�_���6�$so��(��s?�CU���/�L/	v�82KL���j�����&���+�9���</�Fg�m��tx���U��x"����lZ8!��Pf�"T���{X�'f�5��<�|F�A�1��R&�mk�9K'�Ǆ� My�J�s|�?ԡꩀ�'�����ھ�O��Ǟ	��ye���DNix-��e �*f�pt�4X_D���^ۖl_
aӛ�������CwO��v_���X�9�
m�WSBI@�tG8�X*T?ϊx�s��;�v���"�$��dG�$�������8���^�Ui2�4�E�&�ug$yU�Z����Fm�������RR���5�^��4���������L�����'A{lf���n���Y�*���TŤE��ZwV�qޱDW�I����<�}�<y~&�|/I0�IU.߇`����D�0Ob���/�P {���f����ų�RbfZ��5�s���p��o���e�z��}ίˏ�#�ă�WF����O)������xd�m��R�����Mwx�2�?��/� �a��_�=o��O����C%jB����M ۢ�V,ꚍ��
�9 ���D6�{֣�a�خS��f��6����C
>�L4�l'Mir�S2�WC�iF�:�|C��8���"w���Ĳ�,3/^�$�I�� �=!suV�r��A�ȗ����\w�P�\E?z)H�ra�֍Q �>M��U���=�ղ�GW 5�����}�)=�I�m<��.>(�ح6��:�U�*����M~c%m��˨8�ٝ�|��4�Y��P3��L��E`R]����m�:�����^���<����O�� �%���nِ�<`�o��{%�ҁ;�xR�ĝ.i4�����.rI�	d+ �$!��Zu��?ƥ�o���5Z�!��0\��Fo�I1�}�kh�A(ڑ3ݱ�t�x�|ȸ?�ڡ�z�������C�m��T�uU�j� ��Y�7L�,�Q�	� (��~�]�.�a�Bo5�j��#��fŁO��Y����gnY�k`�6��Y��4�Ň\��:~�xf�4�3�G5�'�P���,��;0E�+�x��HLG�R1��b��>s2<"�0�F�a䷣+�
���P)i%�$�2zǪ~��텶n�!�E�*q1���V��%������%S�?L��}���3�xX^�q@Il,0 ����(&㡒H��:%8X�:�_�Q����$�1���Q|�6�f�ӟޯ���:^�ݴ�8���.��Lre�G��V>QZ� ���}��_��^,�Ϻ�${gFվ����h����L��Y)U�XQ��\Ѥ�+r��T[W����qձ?��u�7 s��TO-��O�nA�Z	�cä��0�{��~��PH@��C���������]��}�z��#����X�E�0��,p��V����_���^¸x���q��N9!�&�q���	kX]��O�b�t�F�۟���uN=.0�� (��:
ԟK{o�Iʃu��o���k��]�q=Z��J�p�IbX�2�RTX�9	����6���m��Z�>�A?����qb+�R��kiM���*}�?1�7�=]{�T^���z�95��>����9��sҾ��"��VƬ/I� �eIiQ�����X�<��&��č�J��Q��W��'���Z~�D�i�@��\��2glS7!� �i7�vj�B?�_���4���܏ٹ�fa3���~��W^�T��е.��̎����U�)��ڭ���HbA54>��bV�f�����:J���.�����I�y�d�F:�����v!��
Z���X"	�aD�Q!���N�}�.s0I�b�L���<醗���>N��gep��ou���^)��m��P�%r7�`?{��9Lʮ���|'�1a����*�;�Ӌ�;��S�>��)��8r��j��y�r��6��XȮ�Z-d��d������@�λn��c��y��#@K���"-E�F��_����K�Lu�7M��Q�I0K����.ɶ�պ�ۓ�Ylk���x�/g��L��m��I���v�*J�؆���G��ָ- ���V	*]4[��y	��m⿊c>�����E��l��P����=$H�8���4G�]-��j�hs�&q���D�;�"OaQ~~�P��S뫤u��𷿳DU�'���n����0��Lg=�S��0bd�P~�#G\��z���%���B�"َ푤L^RC/�-EKt���F��-ozL�4A/ϞPT/*A��9w"��`�N�r.��:`}'�+z��Bz�����g�2.��y��F���T�J�/�����ӳ�U��-8D����1 ��3�$K�E���*�HD�����-v�L�f^�ۍ�Ժ�V�CE.�OX �l������s���J�0��n}���ђKo���$���;�WB�W*�>����_��0W�{ul�2`7M������}�%f�ˏ�-�A���R���3�?`$�ۻ<��۪w�|��~-"�m��~������:�66ai�|�"E;٧b����8ʏa�1\;9.�Y-�h��>�|��;广��DCB�֪-b�`�6Fi.�K���c�?m�1�GY`��A|���'�v]۴��P�녺p�
}�m�[iBQ���h���h��(3�1���|����:��(C��
�'��G�G*3�Q��#s�2�ga�o���	��}|
ᡥ�@��CE�c��{�d�b5�WE�~�R6	b��+��uY��f3>��;�:�������YkK�;���_���rR� 8�?��P�&�$³�~���Pxlws����["aB3�X�k������Rn�}�}�d�`�w�ޟ��1�rk+>��XG�)����j�n��-j5r{8D���8�斻��(��~)3T�t.Eu3~KO���4`TR��z�z��)�)��-�M��z<u��*ZR�����Tt��R$e>���N�|xcu���I��T�l�[_��a�$��ۮ�~���Xx��ʗ�Ō�1�x��a�eT<ٮub�X�tҦإxд����әGT=��L��-�WJ���֬:k�e;��e���+��9�X�_�u!I��r`%+����;9��>�c�$��t�A}���<�}��9���3:��(՟���0FX�L���F�flU���V��]G�r��-��s��wz}�Uc�Dn �9JW$٣"4of��������CL�~���3V�eX�����X�������sr���N��t�B��
�2�@Sh���ӿ[���X �Ξ�v
��n�Ð�/ͧ0�'>;V�͇�����Bc܇~�"�U�M�rl��&8��@���Cz0�:D�����R"���[�H(�9�N�r/���8��3�}��������a@>0�Xo"�]�`�),����g؟:�qϋ�� �d����շ�:k�5Ɠ��O沪�*0���W�w�b���
u-x6P�򐤕�b��oC��)��[��T�Q:��5�П'(^�ɮ�S�o�u3]-u�4Ts���D���Ɩ��k?���Ѻ�*�a,mu���0��"�;�/~�d�g��Z��$�ˠ15����� �40�$�bߗ�_拚�Jv�$��ߋgÑ�7����I�1i�xo[#��z==�N�g��^I=�i���K�����2<]�I�T�X���:�X��ǭ���B0/�qв�r���m���A����y���_*(��s�� ����;�?���j�^��';wJO|�R{r��L��(���u$ &}�HX`<���]aY��x?�u�qF�bT�ې4�{+�Nй�wv����h�x���iBI���J�9j4���-#l/���ѫ캍G�:��'�Nv=�y��W��# ��|~��Ђ~F>%݉W\7��;��4񫃋����`e2�F��B�qG���Cswda� )l��Z
[ۨ�/�a)��:��Z�O9�h�gE��q����w�!g�%6��o#�8R_+$]�P����; P�
���D=R�W<S�G�ӟ7�&C�*�VN�3>��}�-bW(+�Il2I���W�`R�4��p�����i>���j��MH�4V֢#@~�!�{��8�&�i3�Ƣ�*�iDW@���yo;3ʜ�8����t��G��Ps�"�,�&��)�%�p~�?3쌌����O�65�sXB�$Y�f������3{�.��,�We:Ⱦ.�tYZL�������7��Q��t���ڊ�p. Ea�7��X���64�U���bT�8��W��ܠ�G�"��ٯ�6��#c&��)0��|Ё�*
��9V��sMD��e�y�uD��i�#��ʄ���Do_�(��xj�	*���/��67�A!�[�52�H[民	۸0X#%����Uk�E'��o����20S�;h��k�G�l�6��]�j8�y���������98�z{� *���Ej�e��V��~��,�j��_\��/� ��#��=�����H]�Q ��	
����k������D�Qu��Ș	F�+��R�I������oY�wE�Ū�b���Y����g��.�04Q�B�t�چ��>���L�myKW�#Z˧���ҭ~j���-A3;
���+�I�e�?�젴#�Ie���������<���~�ur���NԒ7��5�-#��ff���ȦVבݓu�u.~���9��6�t��y��)3@h#�')�}��%F�vOF��Wh��G�=[<T� `�x��ݴ��#�����r$wWһYpTJ��W��)��54w$k|ĩ��ل��<,�S�r��-lP�]�g��(��W�w�j�n������J�L(�����-�����=�կ��5�j�
|_��H��h:9Wo��޳��6�s*5ߵL´gBQ�'+cu����QrG�ah�(�(��ԇ"�7"���
�����S��Rq��������j�e��R��������!�n���$+��Of(�o��`�r�d)c{�$�P�UbZ:6����8b{'��x16�BD�� �B7�����U6�o��x^aBā��O#$���܏T�e����2j]7��� M�w�,��b�y �3cr�g�"��N!�x��b��_S�Ͳ-f��8n��_��G�"������aT���n�Xm)���&�߾���KF�ǡk���p���J�O������ Iva�7�F���}���2�4��ᚶBuQ�ѩ�5�=݉��A>����<��e��hN��n�z����J_c7��2S��:���8�^�Ʊߛ��fl�-G������.�ka2�-�ۛ��4����Z�#lI+8=B����� �@l���2µ��Ö�vߒK	�\�K譃.��\d~��I���kT�
��S(��"y*�V>����G�.I-5�	�$�<�^�i}$Qik��������6^�^�O�܂�9�T��5��K�~�Z�{����c��QRU�<o�}��Uȵ��v��ї5��ӿ+��o)���BF,PUd��4˄%i/N5�_��#n���x�������`�zX�[		ov�����<;U�q��u��3᭘"�D��� �u�	�ҩ1t�R#�����zu1����8��Om����q��gb�9���Z���)�P���Bg�*��.<�B?Nc�����s� �H��zk�(_Y�0�D�em�U�#=�w��S�&W8wW?&R~��= �{D^���[����_�7�1�����$���	"�{�~	!Rmi�1�[C��lI�jֱ{X
e�ag����8�����y�_��޲�~aS�V�9rZ#C�S�]��9���
;������Ɵm}�5GĮ�$�p���H�۵�>X���;��cj�z�r�Ӱ��.�f�{���2'!�~���-ʨ�/��Uc�$��:��V���O� rQ�3�L����(�U#!w�d��t
��������J1�p����Wi�D1��	��ú�*�%�ֲ*2>ڧ�x�a��ԩ���^b���mQA�Ҥ��Q���#}�d�K�<O�1c<9�Q����q�,�Y{B���*&{�v�ͷ9�M�^�ޤd�8w���p���QX#eLvp��ď��Y�.޷7��l�&�-��zT������ca�[#�[�Yl�kq���ȈX^Djf9��6S�{��C��'����m99�X��n��"KJ�0�x��sqe��^h^�*&X��+U���ߩj4In�s�$d��,qpCy���#���i(牀A8��'3���FD���Sx�=(��C˗ ��Y@MQd �����M������-�G���C5�!�B)ٜQ�p�*�n��O����8���Մ5�,�7J���>�	�)����5��z΀_y���m#V��;��q��������A?S���Q��&{k,��6Cr*�Ȑn��"�}��m�D�|�B)�%�Ne|3ja���R� ����p�(�e�U��Jjt��9)�;$J�*�ۘ��]p������4^"�ab�f���z�\L4�R?Q'�=�}����eC$4q�HDz!66�Zv�)!�g$κ" 9x�8�
�gU;�T���]<7�&����j��.���}�C���6�o���+2g%i۷�>VO{Iz�[rI�$k��斕2�=d#�޵���Ct4ܑ�� %J�t�s���됚��x���%xy�l7�ue%�"��8��P]D�t���#`G�"X�v*����^Q��㡦u!��xΔul�
�g�K��Ed�l2��4aP/5��p%����g���Z��z@����	6$��E'���H���u����q���%���k�������G���#�h�zZ૜�n�a�k(��k|��Lm;������q@@`ί����W��h-��-�fF��}1`a���)��VtT
E�0z?��c��`���2ԉ���s����MO���b�$����B�@�%�r7��k���[-�&|�"v*�e����4�*���ow����Cv�3 ��LǙ��泉:2��q�G|����g��G4Sަ�<��==���PE���XPȜ�,B*%;X �&�ɖ�с�Ҍ�l��5�-��C�91��0o����Lݙ��U�|����ɲ
����ʼ�@06qQ�u�=4�'f���^����� F���%U:=`3���1N�F�|�������4+C��4jL��ƹť*5p�O���s}%����J�n�U%�n�v�[ZU�7զ�e�q��>�/�[0S��6�8�Lb�#j4��PX>\N��{Adn742S�MF�����!��s��ຑ�U�9����`�q�5V cNZ�:-�Ѱ["��$��!���E���e�=�AHN�2�<�?�S紦��h�9U���F㱐����]g��"d����it�c�(n&����c����Q�;L%U���uc�s5w�� �]j2�<rJL1+�� X��p�[�7�_PcF_��`�7�Y�XJ��NSFH��M&1�Gv��~K%S=�Z����X0�P�<�Gˀ_�.�O8 ��1	��*opN��I�T��k꾠bάu����s�a�,��Ԉ�6[�F�O<K���A"V7,6���>%\��[������C7?�w+�J4�>F�K*r~ԪOdQ7y5`�~��A�;@��i�F5�uɶ$��,Ѓ�����!�#��kG�4����Pt��kܓ���cD��>\�\G�W�7E�y="�5>^��"7�Ǵ}�eP��Ƣ";		A��{x47!}��Z �<�폕Y�8�g�S�&������ꕼlǢ+� ���W�G�͜�жŤ��>��)��D��yP`�u %����d�B]Q6y�q���kM`ŧ�\�u*�v�S?2z)Iҏ�<k���+ �rf@��
�P�6������{跋�H�K6�1� �%H�`|���c�O9���S�̟|��a��E��*�:uI�{���3��5Ψ�Y������bʼ�,�D1� jS����� +�r�^! ���+�,q���p�6X����D�q��+f��%~� �с�ψ��&��K������W=
����Y?�?��"�!V	n(w��EG���>�D�q�C8}}E������r"T7�X
�=H��3U��O��'��2�7��v[l�!�d1_viN�\7=~��=U��U��|��V4�B���IJZ�J�-=���G�m��{��J���#�Z��@����*�L�M;�Gs����5̌�H���c��^|z���$Q�N,� g[�B3Qyc�?4ߋD�t(�Q�l=Aq��5���D��P)&Rg���2��{�B�x��`�Ę�pB&%�!���,]��nXra;�#�(�{�Z�OQ��9����ql�vr S�N������_^�������w�?.N��~�]�0#P����6և��7�V�(�#I�_������[�p�1C<���a����iS�(Q��D��l?u[>3��Pi:iy��̒�=��݉b��̱�d ��з�(��np����@����L�Ռ��,���!z���T�[�`56�=j{�χh�ɍ�f�0�ݔj\\��h���g��%�r�$e��:��(�]�{L��CD7��5�}��jp�Ű!���҆.��Ќ��Q�w׎�5b��+y�j��� C���b���:� �Z�9��>T
T.2���7�,��""/Hd�kGc�}0΁�sj�B2:1_M(�I'���c�]=��FK[Ӄ+p2�>�1�Ӱ�Z�XZ�C�nr���f���$�B��}�xM ���
?P�;�%�R�Ѕѭ�'kC�����30�@vT3kxbB7�'��(ĖbS{� ��;F�bG��F@p��BRu�Q�u5�S��CT�a�ԁ���}49�dS����U;��a��-(�ѱ�]v�=>țe� C/�F��3-�q�Xk���"ø@}QEyآZ���	��ez�f��C{r��6�^�*����$1=�O��F�3���5�+n����A��ގ������T���~{cz��fl��ƴ����5�3!o�SOY�(�Z�7ϒǢP�?�t�*����	[�ѵ��O_e�3�s{eއ�L'��+��oB����,�6:K�&�W�ďp�ĥ�2h���S���&g��:h��|��H�-�M�B�6��17H�$�9&�@�8gls������[XybvJ8��xB�_<�ʍj�HF#�WR�QQY^%�u�ڹ��ٻ��;�'�ݑ�� �� ���0Ɩ�i��xp�d�fے ��$₂���Oj�����q���J�
�.��������>�$�n�R�,b����鷻-��f�e��� 5�����7ۋ��K�C �cv�n�M~�Ԟ�3��ӝ�n�BtIŊ򒪗)Ci�>T9��ʡ���"���H���@�4�W`�f~KD�����7b�G��?�#��i���dwO��؅�!/83���ϔjO���g���Z�\Y_o�������.'쳠X��ķ�#����s���<{�'�-I_ �1��c�q�gI��n�m�R�:��MYks���`��ymM�Έ	ۢ2�qI&1U�[�k]�OI"�w'HK�y�(&F/$�[/�±Hg�X��_PA���*��F��)(����\�H���߫%�h��ま�|x��>�v>����H�] �)lP���P����Ǟ��w~��4s�I;�� L)3L!��UU���v|u�����8 ������>&U�`�jNQ�C6z�\��*>4��dxh��m��6ԣFNN���{$Z���0�hJ+B���tZ�b��탺R��^��3�!��b�LW�����\�e��d����G��f�*���>P��5{��k$+N=�u���fc3΋��QL2�����Os`�./�g��+��X��ċ#z��f�{�3y��Q�v��a�Oe:�w0^����tA��GW�!���;��I�}�T9Ga���N��*�������i��!��y�˩�e0\���R,�X	�D��q��?b�)/_fj�(��/��i�����\3��r��c�'�J�d_a1g�fL��;yz��	Зk86
9�$Y�L�n�NѶ�����B��t�u�T���J����A��/V�3��	���UI�@Ê�i����P�H?��kSp��J�?�W������Q#]0r`�!X ��!N1�jS�%Z��[��A=�$R��?�Bn�K6�m7�kBF%�3�ɼ4r����:}���2�:N�in9:�oP�Mb�%���i��q;�4ju E�\��)���U��X0��(٘��A�G�o�|!�+}��̓}��	���{��	֒�v��Ī\G9r��w^ ����&��i�����+o� �{�;��A8��7x���67C���Ll�/�[w�=���Alj��aD�Fa�}�	x�VFm�_�'��ǰYO��ڥ�"��� iN��U�6�˘���JHྀFY�HEMD�}���ygo�fS�4a.��O�c���G���X���K��=;d9�C��i��d|�<�<��]'�]=�W���:�+`���y!F���h"�#���x򸸎�����l���g���G�5ܕ/(Od��ך$�d%4l#j�;���D\H������)M���_ڵP-7Sӂ���H7QaDYD����Q/k ����C�5�kvbb�=n�y����r&m:�/�IX�H�+a�����wQ���0@��k�N�x�+F�7vU�Ɗڧp�_����F�n�"U���iL�5���A�r(����*�k_��6\ob9�����df��YhI�f=B)��]3����`k�!x��g�����2L~�,��*$��"�E���|{9eZz����l����|(!_��QV�����mV��H�\c_��q����>�SzpאI��0�d�������:tLe�ӄ�f�i4�#��I�Y�M��>�������M\����)9�9݌���I�b��[�/5�:|c��+̊�q��~�5~�V!�M�.bź��B�i��x�!��#��$�,:�������7�A�!y�'n�O���̱��[>�KfA5�(0-�j呄6s��\�.�f�k�5gԿ^`���ۇk	�7(
�ǕA��uQ�C)Z<덲�M�����_N������l���oC��N0M�p 7�ՙ���:��z�|ˋ�mV��s5���
��qr˨�GXc��;��p��t�bÈ
R��c�P����?�Z�I����;'/��,�Oc�ց�d�~.G�C+	��Ѯ��`�g&����*!�1nС��*��=���k��I�ܪ��][]b��2��2���]���K�_I�)��}-*���96���s��pQ�VY�Ll�se�#�0���X-2�K�/BG�|7�}�&�D|�X�@�>N�mꙐ��w�1�ǿ�(^��w�NA  X���JJFs��",z��-k]@��/d�Dm����#�5���$f�a��G��@LQX=lu��B�Ȭ�6x��,ٚ0�"�aH�� �tTx�u�(rn��p*�)s�������{�����U��J������c=��Ԃ9�d��d+�F�u8�3�~C5�-IܥO'Q�Ӆ2��Gk�=�)hg��Tͣ���5'�z�����G��Uf����yxf�܃h�+o|佡��$�H%�ԩh�����m�,D�D)�_e\yC��}^j{�	�y/�4%��w�$-2��,I�E�~b�g[��gۺ�+��G[�} �a5aE��Nu{K��|%�|ZL:B���ro��+��'�E���	R8�(V�#I����0{�}���������f���^����%������˩c>�IFce��M<y���۠�Y�;���Nq�#�����=�N�u����`B��o��vp��E�J_E˞ݦ��ɂ�-���/�-�"�����`Tǅi{����FԊ�i�4ĉ�a� �|���ń�����`>~5�ǆo!��M�؅�9�s!�Q�� �w�Nz6]��2ĩ�,F��Wf���*�E�ʑ8��~�Z��>9U�3'�X�$�4�?E׏Ag����aN ��o����g=w������&�x���z0��o��]�OY}5��r���50'�)��=(:$�2�<���m�vWƅWt(ϑӫʠpYéJղ���y��x'4�	�q߃U~���}�"藂��F��~-�R/�_�ԃ��EԳ�u5˝�!}���r�P��űK�w��H5��<��u��\o��f�A9�b&�t�h�+t拿��s�j�n �o�8��%�6T³�/�e2���C��Uoy�-w��m��pt�V�kȖEn�'�%����4��:=N�)��A<�[X���,����Ul(�n:�a)�1A�5�$�u�ٰv`����]ߐyC��*jݝy�Vh���U�Š�9��^p9r�A)V6N�c	�U�
���o?V,q{`+�zQ�:D�jnԛ�xވ=�쬱�S���h�*�����$Eq�$�j� �f����e��΢ͤ1h��¢Wu��첂+;NE~��j�e)�#����j��h��$�d�(� ��h5[�W���L�D4�L�{%����6��ctLڝ#�A�]�H�<�r��6��2������2��o����?3��d/��f�*��
��W0Q��9���G~�Z����(���j%���D�ccףOa�QC��u�{�!g��m��A���p��]�g#��Iw�T�S-E���^��O�}�^���ǽc���CL;��_�Ӏ�d������f����[�����1N��� �y��!���r�P��Ҧ�y��������U�����LV	���L3�3���t��K�4S�UU �)q�({yq�r'�wV�;���ZΌQ�`!�:�s]�hw<!�h�*j���7t28y/[��F�.˱�/����|Ě���m�б�����?�����¹*XqC�fj��!��6��1|����p���Ċ͈���=d铪_;�#-

ҝ|�ы���n�u;5Y�ؔ�Ӱ��4	�c�opL�z�ip���x���UC�c����oy���{��h�0f@�9>.���ڰ��C?�"U���4Ηw�$�~'�r�A�w)�|���O���� -�M��A�
[(�9�M�0j��+�a� �jd߷^�ٌqL�l̤�v.������k3�B���uD,V�Kz8<�1}0�d܀�)���c��Y��-�p�0�H9���Fy4��\��G'���,GBR/��&� ���p-��SE�P@7<Bh�S��õ�S%�-��P���Af���	4l�)q �ҧ�4�,R�?�
������)щ8y����PѶ8zX�x]��Xۊ3�/�ۡ�ܮ/8΃_��X�����%;Nr@=��g�X ��{��*Zb�m��W�-k��4^v�s�=�<S��!��Z���Ȟ���KwO}�/��@�SFq��;���~y��*W-��0Y�jg���p�ƫ����Rx��񍾹|B�.�PW4!���6�d�M�C6�^��G�����^���b���	1��[�ՠ";�˅��nI�`���JI��9��7@�8[�c�%S� ��� ��q��.<K��m,MӲ`j�R�ǃx'^[5�"D�c���[l��0��4S�ī�^xɞ���/���w8v�w��l*%���\�����PC.r�x���0�ļ��E�,Im�a�;��jvf���p} X��o��.<�5em`�Vt>����y�3��Wv	�S(���(P9��qQ3�+���˔�.r����l���w R=3�Ӆ��]Gr
��{��������+�dP�������j��dpA�yGfN���ޏ�d���*!�平l5��öar;�����[W@��h���{��M3�״B�[K�*$B�F�xu�A��#�����۩J��)� v ")�����f�5�����۪n��8xD�*�+�vX���a�e��gu�p[���
��I��g���.�O�6�?���D�� ��9�@]�Ӭu!�.�6[cU���g�X����~���&qĞg��k�zD/	�G"�r2���"�j������)0��L��چWJ�ꮀu�vX�<We8,��Z��F���)z�fR(�zZuQ0�����F�M�3�Ƅ|3Ӂi��ߗ�hޢ� �o$�厦'-_�}�ʳ��nU����1/ɽ@�&��x�=^����0��K���?�`�-�C^�O:C�(�Fޛ ���]�Oٴ�a���3�>��5���~�e��|"�iz�;Ӵ(��kg�jK�T�ia,Hki�鬂��M7�d�̞����6�� ��/ԣYU�P�6�*�:�AîU�;�9E��Q�­l;�	x"u�/ ��L��y�a4�(�{��&B���k���lj���U��F�ރ}k-T��]Y�hlB��-d�B��TW%�O�zN��u?��9GQ�`������sDx
k����w�Х[`�msZA��@���_�#�T�[d%�0:��:n�3_.���s,`���965��b��Xѧ�a$��\��@'� ܑb�,�"�cpO���R�R��Ÿ��+P�}$VtЙHN���Q�{K�3�ɗ���/��XA)�9&� i���<b̂�4�58�c�F�Q
��X���i���M�ͺ%ݛlt</J{梼�y��
��~�e�Ǵ�@LX1T�;�l��!�v�[��ً�o�l�Hq��e�soLP���B�Y
��reY�}a�f����."�;�
<�'�M��� <��>��*J��5���������u��	�"���~)�,ߝt��������շ�|k�ؕ���e���4u=�����\5U�`��W�x1߮BR[q�z~��g{���ɜ=�!��m�#N��
~sŻ'�(K�(��W��`�1��]������h���غ�Q/W��{c�ZD����b&^P_�.8{�{��c�c�I���F�����-���cn�^�,�a�/��9��2�3_��r(�Y�3��cC]��M�S#��p��C�K��*XV�u�{���*�o%�s��c���F���/�w��꺥�uJ�!"�Q�?Q$���F�n����Fi|���OҌ���mzB޲h��R�����Y#���/m���Q�1�#g��t��ޜ\EX��o��g�0ן�3D���2�]�\��.�~Nk�c�{H���x��4���V��|����5y�f� B�X8]�:�#�	+�j��k1�\�mX��j ��dB�������pgג�-�cKd9"ƹ�D��!:�=��+��)o�?�X)��{�t�����K�ۮK[DP~1��H��6���D^o�5ׄ`�I�At��=A��g��p8���y�\���)�Fo�ﰻsQɓf��7o��u�#e��;<a�`,��&z`���C�sk	U�$�E�'�w�;ڳ��$����I�d�Y�&�&�1�*����dj1��L�,�,t6/Ⰹ�8iH�2d �«V"sg��ƏT���N��%�Aĕ��>���aj+N<~���Lu���5���8�s�Ze9R(�����˗6"}9��?��Z�hʣz��-Lg�g\z�"���b���Ĭ�h��{��t���qm�Y���o���%��UYB�P]$ҷq����S�d�D���5)^XJ�\G�D��V������|�a���أ)�-��@������%�W��&�:��~B��Uo��LK��^#
�X���LJ��rT�l��{6�e�%��������\�Z�]Q@��Q0@��^L[����B0X��R��EI� �](9��%3�-��ڼض���A��2���լ䬓�zP��,�Ԉ� ���t��S���w�;7����_<י��W��b���Z9<տ���K�5F�Y��d�TZ�o�A�����.��?���g�x#SdFS�t��+�✴�#&�t�Y�x<���N*i�t� �S���ZX���.���Ggj!}��XC��L54��*n�P"
��HS(���U�jk����?�aB�%6�͚���.;bGǹ��H�U�5��3���9pե�]�������ĥ�NzFq�5[��v�U�g����~w�{wEC����"J�2!�,{�����n�T6\?��!�9.ߎ��b�e߂f���(�t���>_;2��%�;9G�R�����imz`Y 
���W8c��D	��bJV�&OM�Q4�)�����J����L�M��%�4��~:���D+wg�*`㕬�P]uN����R���[�W��`��@�P��P���اB�ݵL�Y%^�ޠ⢑�=+D�,O����J7儘 �2�z�^-�El~�o&9�*vj#3���]�7rZw�,EQWbVZ�[TS���}cu. �JSg�7R_����f7u+z��u9X Ӽ~V�.@�� �� �8dG����l�!��ի%����]%D!�v��T��&� D����%~���2/`ըrO#��u!(�����9�!��d!xn�7����ܜ���=�T��V���]E��~kn�[3�'B��L�q�DF�w'|%�A:/���X<�l����;(����l#7`�s��<�g����^t�\El��[k�a�~�w?���v�t�M�7cC��6w�bz!��X3������WĖf�ܟ�gP��������LFJu��C���"M�*I�@����U`����S����|i�C��P�W��Y��3i(��$��Ռ}�?X��@K%�=��-�߬�#:{�2Y��	�Y��~��X��o� vW1eֆy�D��/�n���"'yJ�lS�ղ�~Z�%�ݳH*&�N��r�Ų49:�e�M/��[����+S�"i9x�5�5��.�����Lq_J��L��� �"��:�T��r㘙M| ���aAMO�s�TTC��#sg��������f�ʨ
��_eMM��(b�/{�(����١����㤯��Э�ǎ�z�>P�f���[�G.
1�D0����
��>*�|Vqi������Lˇ�hZKZڨ@-yj�n�O����0&Xtk�l��͡��Ty)s�u�����"�l".�s���O�j�����3S�Z�j�C�.�V0�"~�_�r7[�q_}<�ive��!:�5�ሤ;�f1��Z"��nΓ;��7L�w,��^#�K��2^:�鋥�O.pl:&�9�v�I��F}Пn:0̲�Fmrn�I�/�N
T�u/��ϝ߿c���H�s�'x�Nb�0zzi���>.|Cl\�&��]%>Э9x�'ȔTŬ#Q�莲�����(��;���x�FT�>�$�����士�W%d���������X���,�m�ݍJ�"a}��t�!�`+�ڡ����Y$�?ܲ������*v|9�f_�s��V]��J��nd��%忹;�Db%���[����/eOӁ��L���C���&M��d͛�/Ǣ5������32g~��z���!���%��g1~�,��y0�w���:�.4�L0��n�����R�3�q������+�BI�rP+����%��oeO,2����\���m��,��L�ql��ۆ�Z��ԟL�b��^��ՌL
��YaǄvv'�o��0�_�^�i
����|v<b��q�ZMޖ��6.G�Hɴ�����e�~��V0��藜y[V,k8�:���y�YHP%˿5��5���odqf"�a�HS�I"[�2-����D��V���klM�LA�B��eI6e�}��_!�1qA)P�x��R
M3Y�*j�{閾�>�
�z����\�i����8��Q�x�K8oc�s��n�&Gؗ�%��\����8�}��o��f�M��l��3肸��~�*5�L����;C�G�)��z��.�8W��Y؍m��XY���S��UV��` F^N�kGK��$3.8z+V+HeS����}kak����,3�Ζ/Pt�=����C��eU����l�J��MࠝC	_ŗ�z�����
��^�\�B��>��+�e]X���f�l?$��J`#�NC���0�ބ�F��|z劰��|ix4XX A�(o�4�둉�/����;ҏe���M��~��Z��g� _��.ǣ\ۤ"״ɷ�`�U�E`�i2b���xW�V���N��ɧ��Fh���|�7e���娉�8���B�JB[qn�#�+ B&�~G�5k�@�3 �҃%���G#.)* �����Ex�:����p���4�n��8?fI�D>p�77���	éёpN���\xkV9���q�i���+$��]�n$�;u�*/*Ա�>�5@l4��iL���Bf�=��}BR���xc�_A���&�ʐ$��k��aV?ڱh�\i]u�\��I!Z��O}�H�D�hS����ry� �����Bb�"Y���]0J��~U~Х�^��[T�U����F?_��Jo�P���]�Q�M���� �3�¤�y��2��ի0����XM����
ߗ�>�c4�K���ߤ�/%խ�#�����)�\����,���9|~���w�K��`��i���_��,slC��]�n���i�1�#+�)\:I���>�(�cbK<��(���8�Z������j�V�5?���躅%�!Q��������%�c�H���H�� xwr0s�������1j��ȴ-Q�i^��S�2>���l�����
����r~�26.�e����3�DńXW��Dƿ�"Y�ڈ�L����z{�c���Ȃ�0��u>h,Q�>ko�r8��X�.��=�`FEQ�h�UJl�0��<�~P�jh����L����Mp�\O����;f)i[�o�#�PV�͠�9�}o�_������_���$"=��:6�<���/=�K�?����@���xZ��g��� �hq�4���x�$lTɲ�B�;��}#��%bʔB�l�Yi�(�0��tL�������^[5��IT���(u�8÷7gKzu�|��a�Ī1f�(WNr��'\�����NIii�����lS��|y�E�or�@����rg����nC�.G���\=����"�����"�n�G��B��)�'}NИ���P��,�x�H��ݰ��=+�"��n�煮���~Z��>*�is�X��M2	��N�g�ڤ�L��$���c�vaω�Y^������G$�h�=|�1��=�0(uM�Qm����;�Y���K���\yY�k1���d�c���E�B���=v���)�u�v��>z9^�$���H��r�M~]�f��2l��'W��>H+2�G�l�x����4����"�Ǡ�x��`y��-���4��]r�CT��0�F�
��0��³Z׋�;+S}@��B%��չ/���=	�<��B��OyΈT�KQ�v��ybtk�ϼ�@��.o�'1&� ��Q��p�Ը��36���7���c�P���X�}���r�C� Kݎ�"��Fs���?���Z�|zw�N܄5�	7���8-4�xSߥ�;�!-�x���c�`���FA;�����%�*7A��xA��LC����}�05Ԣ5z�hȀ��u�&���86�wB�2I�A���6��ON\����2��t�k�\N2�;Z��\�3�Hcb;h6x��&�s��YQ�)v�E,cダQ��K&��]U�Q�MJF�Rߎ<B:��_���o"��_
yz@t'\ѣ�"�**��W��|�zqu�<E��s��)�q�m(�$ӞT���{�_����:�4��y7�$�Ho��ܠf[�:�0��"���� ?�ۙ3'qƟ���N�R������Ka;��Qm�r�1x���+o�C&"�+)h�P8r8#4p�̉��w��Zzd4�<9��Q��g���~M$MO��ݪ@�� ����ͯ����5-O� -��� >f��t,#L	B��Ga��Ւ��i6�]p�C6�R����b
���&�<[b���P}�Y�F��ē�q� g6�������F���OV�S9BRV����V��%�#��,�>�ѓ^�+�OI�:�6z��x��~q̞�CŃ�f���k�nY��	0{d���CkL�=TΨ4i�0E
��P�]�єJ�l#-��V/�Ε;o�Q�,U_��`he�S���"�^k}���X�JOP��d��F��CP��]h�@J��JQѣK[��ʆ��(K�Ǐ~��FoB�Y꽫s&�q⬵����o���Y�<z�hZ��dj=�[�FJ�(�`�Z�I�ԥ�a��:�����|�b��D�[�M��i����n��GF}	;���#��c	�;`^���.w!���w�ɇ�O[�oyP]����M�uڝ��:"a�w�Lq8���"�#�`T�i�Oڭ��ˣ?U��}d�q���h[��+[��F|]a��3źk�֑�?�HM�!��I���AT����1�Zl����1@�Tj> M��%��2���9��ݟ�`޻�!��n��_~H�,x�_ZVw�OR�?W�X_�&�;� 7���_�� |�}Ď�_�4�݅�-�#k?$�3��������T��q�%���ᴚ�fTesiK.�r��I;�Ra߈���Jr$
� �{.��Қ9��H �Q��ϓv��$�4r�8f�l����� 'U@#G]6�T!E��-+����Ki� %U>bi�����j���(l#�ϣ<$�>�_��/p��Gڀd探�����c��̗Y�,0
��w���)���!��Q��P'�
�Ⱥ���������l��D��v�А��pNB�{�^W%���
��bo��Z�H&�J2�%�4ʤ$���w�uT��X� ���~�V`ɞ����S5j�W��F��^�	{�W:�$M�b�@���	��=ֵ���۱mw�l�)����*Y"�뽹+�w���A}�y�i+k�����:x�4���*��!�����8K#u1���Z�Z��J�Bַy�0)\���^箨m,�,�l�����lnuHR���ÿ-��Ct���g���B�
4��y�}��SoF��GJ/%�;DB ���6�t�E[v:�?^�|���"�rWW<�vNCj�!IhC�F�`�s*�$إ�qV���Ƃ�>{�(�4�i���5�Æ�/L2�¨d(�����ĺvM��������n���MJ0�'Dm[�D��R缙��C0�3@rW���c����]��fb\ޜ*�!U(��&!��"x��N��h�ȧ�F�.̄���C�W~��'��H�������u�3 F��G��3�?���	�fϮ/Zc��χ�$����:+�D��r|oTu?�	 �(�%���R����: ����cL
��#�@��F��3Ac�l����Ҩ��������������7�C19q����?�X�^�S��bxb�Q��(
k����G�Y���oa'�����]"	f~.�D�}>JA�A�$��G:�n =.!�L2t�%�3Ok�q���y#�Mm��iG!�+\�N�gf�Sc����&ծ��6.�� I?ӆ4��%/�ς>���H��B�Y�����6U�h@���L�|����S)��݄���ҍ@xdt�ޙ� �U��c|!D�~쑡�v��Jhp��~ ��e�cx�$��!<�:MbL*.�CMK^��3F]��|#�%`�z@�V���>����@�L�O�`����[]����Z���y�~zeM���E?��#�	�˭��T�z�e����4��;�Aō�4�C_�^�K�-��\~8��c��Iɜ�M��o�o�xOD�1���g#'7����I�/,���%���U�=�#l7�����g�\XJ �3ϐgm����a4�.��9�>Jm��	t�����~���:��5��{�?}��L���q����`5�(��%Ti2�kR`�ބ�9����6�Z���|�k{�#��i�<ǻǚ�yڪ{C��k�b�r�I�//�<�@	�hq�s������
�p~; U	\�w��e�6B@�"�m�J>?c(��2��x�78�{F�g
��N�m.]:�!���oNC�\���_�#`^�	�iII��mw{�#V_�E�;��'��$P`V4�c�D%c<9(�f�M�Pv��+��,�TϮל4��B#�_D���j�U�1v��#�7�h"+���β&D�BǽQ>^Z�~EU�q���u��S �+�y�mNz��D�.3���I���xZ[�d�1�J�f�Ư8ғ�x������F��Ʒ��|��,s��P�ȧ`oǞ�J�+ܕj8[L��:[V��5�1h��B�9������ X>���X�T�
zt��'�y�EF��B	��:*��� k�S�Cz5U^�Q]��n�H��=^��ʼྼ`�p_��HE��[n�֡������d���m�7�V�=��W~F�솜�/'`�L�=��7dY"����[g�qv)=�Zdm�.�N�	���v��G��� ����0D�� �ۨ�l'��F3�V/*�t����S���|��bBf7�a�=��w*m�ڬ���(ټ�,�B�x����ބ�{(��4;yK�u~�Q<�@��^��:��EO0V{ʖP��)�`��Ԡ�pd�%��D}l��¦}�ِ_�J�C-B��b��VeO���{S��Ȕt���w���d'@䌖;�� \g���Y�F�!u��Cx{Et���;e�-uc��ՊǷ��b���w������Yn]:���#rw�zHیƼ���_42g�t��O�p`j�I��������L97,  V��ƞ������kO��]&�=9O�/�88b�����7gCk�6a,��$2?D�n��F����gx�&ޅ���7���*b7�q�����6����KL$v�F��s��\������/�1���o�WC�U{�13�o����p�o�6����ٿ�����5;ʟ[r^ �ad׸��@ur �*CI�S�����mI�Z���g��Ykm�5
^���_�!�ї }�Xd"���
:�.'1��D��o~OK�B���EQ.3���LFt�V�s_��bb-��䐚�5�MpRM�3�s�? 9�n�Ҩ���������i��y�_�G��x���ݍ�.�����Bq�������<��{���6��O\�H�S���gTXD�����׏i��Jp��a>BF��˺Q��ɓ��\���t[�wZH��ڴ�do�t��z# ŸC��w/���y�����U�k[s[�\J��W�oa�C��	�1ԕ�s1H�wŘǔ��A���7"xɝܡj��?N�e�g�q���@�U'�؊y]�2M^��'��T�ކ/�XX��I����1u[�fK�z]	,P��i����x�$&���V�������[���A�I���2rXo���Ho�4b�B����F���~Hŵ���GB�J�j�1O3 �����.V���MkV2Y�UJ8�ӻ���q���%ko�
���3\,E_[��/���p�`	#E�S|l�a�W��C�I=�m�_0��Ԁ٤R��~��b��h��HwߦAf�0���8� �өF7j�?�$p��w滬�Z��T����Ů��=�A�*�(�����M 0T�xx�1C|P�C��7)���Վ�g H�"��S�{uT����� �|<H
�ć'[Z2}#u0�tKqi��P�.�]"/��ժR}/��$�B�Y���2��دra��"i���9�d]�|�e�ڛ�f+m�e,аw�R?P�s�C,�2@ѦSo��	�*
y���Qĉ�zv��p��ÏO`��.��n��Q���<���g���'�n�9D�v#C%t�G#��&���o�&Y��d�B������3�!5JC��v����bEg�۩��X��wzLa�=�X(Y� 5����pa]�	t�O���$�����ʾ�.K�����!�B�qz;=�=���I2�j���	�
[�2��*j���/�fu�w6Pp���Ku���*�Z�s×�[ �0�J�tt�W5����-|���"#u��qoЭ���Rf����  �xIs���70�����?�)Zp�t��᥍����UC?rX3ݯ�3}n������,����I���]rKIo�C�0ʼus�_���Ֆ<jIu�g��k1
�J3lh��S�n����O�QẸz�W�~�b�ba\<�`���U�;������S�-���F�$UQU��5��m�������!^O��PN�����Z�T0N�%d��4�����
���Ez#�' ~yCO�&3uZkt�̞c��z��b�GA�}�7�y��:���G��7��C�imu!Y���a��x��4@��inQ)x�&��!2�NX��d�-�/�</��a��*��WqJ��?��v�������7�t6[Cm��\����& b��I�� �D�ų��f��h����â"@5b�T9V-�ZU �%�|"���3Q+�ޠG�W��\�S(�/e�FQI�_PT�V����� �H��7�!L��6��x�����R��cv�`�,�u�I�>?�X�(v��%Α���]��Xe�d`;�i?Z���gҺ^�1�KIʈPŠNT��J�`�ke��?��M5b��5�<M&؊z>k<�)���XK%[(����+<��wm��pH�[͚r�%h��"��q�~b!��pP�ѡ���C/��?燶�� |�3P�ؤ.O�~Z�&���?���SV�sfg^@��4u�W_&��Gʪf� ��Ξ�P����i�Y�Ţ ��.4'H�a�$���m;�x=�'n�s3{�iL�=I�$.bбH�!&<��ƺ:�,^��.!�*F�%0�t���h0\�x���2yWr1�V����Jr3!���89����Eh����ׁP��u-*�����T3'9,Z�+�n`d2~Pϡ��_ܐ�ش�Qvm���}`��͋��*�������J�@�;Xo�&��yW'"��6)u�0ن�J]��w÷��f�]�7v:��E���v����
�8����յ�w�j'��$m���-�sG�*!m��ih��!������xZZ/B*%ڥΰ]6<q}�L�R� �J@�rhk�v�ڇ{]�p�p�J5��(��[]O��ih��fodF�ǣ�9��τ��� [�D1�d���8D{E�Bx�S�X���O#4f"��7����R��B.F��+-����p�;��+^n�"#m�I,H?1&P��z�ZBr�63w�x���v*�x���I�l�Ry>ɴB	�iE���(GFpkH�G����Wa�+��|�Y"@K_������Dg�)R�H��@2�۽:^�Rd�e*��}��lw&Ȱ]���S[������`���5��n?�Mu����5fZR�"�����FL����)�v��"���H�<l5�Z��ŬV�_FeC���1X��z�ٛ�OI�t�w��< �n|�U��}W8�|ݼ鳧�̡oC�I�N�0�)`�c��L/��w6Sl��|�� �ؤ�{FK�:��W�$c\yPp�O�/ٙ:	h~烦���noa^B�����z��1e3݄�w1��@n5�* ��rG�f������EG�2-��j��Z���	�������x�\%ٴ֔|���.��"z+�}F>{�e�\L���SO�X��~!��g��P�<V�̃Q1�@R#m�P��B�0i�:t2Q��-�l�_~2Tb�~R��~V3��N�CC������^4����ez�x�J&�j�l�#~a#����z�_T�5Ef�p��#�C{�=�$��M���W�D��錅}o~5������ȉs�y� �(�F�2�����>���W�@�u��9��5�GO=į���&Hcw���Q��W��~jK;d�w+2qڝ�d	�"� ~[���O��V±�*�,a��^ͻ��g��v�y����s�t�A�/�wZ5
(��
�%ͩ���N�\$Y�b�0K�t����~ �h�W�����/x,�H��j��Ia����ـ:P���a������ �*�~q�4@J�kR��+d&��߂'�	��TƊ�uZ�#�;��T����g�� y���;�ʷ�jy>�FI�rh�<�B���d��/ޞ�)�V4���� �!Cw ;,�U|E���0��$�s���x���h;�Ó0{�t:���?)�x�R��g'�1D9K�1��_��X�4�`.��ygk�;k��B
����ޯ<���h�z	I��;3Y?�{���͖d��[�D�B���V@���m4ߕQڣ��T���Ĭ��� $u�>'Ġ�t%���Q3-�H��F&�V8�
\�!r�2W3���#SHhb�d�KA5�Pp���2縧 �j����=i*4i5���b��	������Խ}^e�ja|��<^��Z=\����
a��!Yn^������Q����m�HpG;��ƥEr��~1���ֺ������.�is�-���$,�6��D��id��SC��QtB���<E?GJ9�~hWh<�qLY�Zv&	�A�d��u1�����O��x������$;=�!d�'�u��M�v��T��x��Y�#�,65I1Y\��Kվ���ѓH�O%��RӾ3����H�;,JdQٿ6��Ѧ�CzU��\�Pb�۩Z�a�A*�`�:��
�Q��䰙#Z����F�J��F��2�g\n/&t0i-v�S�P���0�U�� V&66~������U^N��eL�1Sݺ��ɝ�!��'H!��q�c��W�n3�JܡO�$S����Ŵ�Igg8W�,�7� �n5�W�զ�9�� `�#Ө9&����n���m�/���aa9�� ���k-��Q�ܻ�����n�ZѾ�a���P���wZ���'~�)�G�s����q9��E��2cĠ�ޞ~��i�ԝ���.�0�{��s
�&0o�D������þ��S����U��E	����}�tC�V���3�Nϖ�F��EL.�	�6� ���r�R�^U-x����.�tr�⾂�]/~������G'ig���W�UH���eU���t��{�K�S�C7���\O.�S����^o0�����9?%���g\�� ��q�Fւ�W����΄�}��b����[R�]�nVU�H���E����`q8���ӈ���Mi��k$����ͩ�K����5�gu�M��˩�� r�">PC�-u�}Y�Z����
|Lk�+L�kV����:���58�����k�����ޟHVf�s,�T#��cG��p8X�q��!���㟫��c6r��o�-`��������d�=���Jb+xG�pZKl��R�*PQ�=��{^Z}�[-S_C�b����"���RJ߀��J*<���$'f���\N��nB���>cJQ#��H~x��g�H*��Mj�O:�щU3Qk4�D�(o@TW�n���j�uL:M>�ڮu���+��$�@����`dع!����%M�Ǳ���in���Mh��G��k.y��6�Ρ÷���@��qr�/|7��j͡=ѷ;�����gd�Kv���Q�ƣ�i���ʓ�N����c�+�r8Ǻ{3��?g^�5��g�*��68��]21��W U��U�������A3�E�!��+�8}(%�8#�#�,�ݭt�Ӻ=40���{��&[a4�Z:(>����5�v}��_J�O��e��K$��ݕ��OR���:{��^���W����:��Ώܻ*�B,|���ӎ�wY���J��������3E��$�G���ܼqf�ߙ�	�P䯠�n�7Sn�[n����)3u���l�v�^��h��D̏��S�/�^�\��ɚq���N�b��e�,�}=}٬�,]��v�ͭ�׹tk/Mtã"��o������U�AA�؇J�~�:��[R���x���1��Z��ގ�E��@�u�D�����i���i�]p�.�|UqKajb��ށ�,�	Dކ�>Cg8c��\0i�i鎮p/<"ɸÎң����S&W	��zx� ��@8�{���Xu���B+�,�׎��f���酗�'	}�p=dZn����Q��� GR[�"�� v`����Q���}�6�Z�mE�j������HӪMq�u��U�>�;9i9����m�A��>��?��n�E!�	���k��ä�Ŀ,ӱ�oVf�&R=�.}!Ψǘuo2�hZN{����
*�5	m�C��K�$)�ģ��O�؝���<����qU�*ߌ2QI1xw�$�L� 12�z���a�ٖ�Ǔ��J�u�e,m���N&�e�!l���[ΰ�`�R%�>�S�X1^ۦ��cV4$?G-�_r�+�6��O#�F����W3^������
���G����TAܶo��Y�� �C�Ηz���}�
hհ�6>2��f��䞬�]6�`˗���w(`9j�͇آ�;Z_������F+��m��ݳ�����LB����$��,�Ǝ�hB� ZEh���\�!.vDM��&�g���Bw�M9"3�Kk}H��I퓆;B�G8��y�]LvO�me��9.  "�l��}��Z]1Kq|��!��r-�8��r��d��f��'�d���#`	�ƣ�8���KM7g;��$X�Km@b�&a��,Js�.c0�γh�{��sM.�H������ʧ��8����l��0��h�<l��&&����7�%p����r�σ
�����}����k�8`�b6t];��xf�me��^[�B�M�~
I��Y(�T����z�;[��~�lck�cF���Q���#X���)`��`<��s?�����A��&���G��U�ɮb"W�}(�|����>���S��fqc�m�Qy�7��X�ӳ=rk?,���(���kE�:�.��0hmDn.;����/�Z��2�SD�^g������Q�v���_8�B�ɘ��� V�.cԙ�-9�A��Z�*�` ��P?H�ױ�����m"�N�9� `Z��l����S��������pa,�f�&{�����xa�u���E�A�FI�ߧ�0��6�ᱹ��V������7�E���./<��Q)@���o��T�������3KH�H^(�%(���v���C3�0���Z^&i{�J+!?�s�^�P��Ƹo�N�C~�P�ō5�����:�L�٨��T���IԳ�w��5|�ER������"	�y�e�ڐD�7�n!/��-nt'-׶�6���9A���U�CG�!6��[�핹4֕e�]/rּ��tH�E&nFd@�XD #Ҟs�N�ȴ=g�)Yu�'���dT� �}�v��;���Z2�g��)��p�wp�@e���*��@A@���J���NЁ߱�g����_ygٗ:�W��ȠrE��l:�qJ֏���X�Hד�L@͂
�[bo�|'(vu��Ԗ!̜CxK�͝E�&��cD�%@��v�P���\LT-���F�-���r!�o�
�~J���K�����K
e�3���
�O͉�:e�e?�r�oy��b�L�y%}�ľ�@J"T�nRo��*4*�&�K���[�h�ʖ�*�s��$�$�����s�%�m*��/�z��S�%B���/��(�w
@��|�D4|)�i�p�>��ځ��������&<��z�ͬ���U��N`-�a�Xo�9��a�w+���q�����J��zy��b[-ul�,ݡ!7D�:����V�:�2z���0�q p+,ݰ�z�܆�i"��!�n��%�V.��B����T�i��H�QߋG	�h��3���r��[��v��_ސĻ?�~�pA�$�����2`e)92+U���X]=,�Xfo��-��9z��E�� �z��\|#�btm�e����R�����j�%�t�iNJ��)b��FZjs��oY�����O�m ��	�A�W%	�H)���ͦ��h]i	�<x+��8a�h/�4�k�龡�Rqf>�@-�Rn��e���V	���k�{��}��d���X���Έ�6z���_FG�qz#y���,1%��d��R_D��EÄ��b}^�z��a\ϩd@}���2�����g��7�3�z��d����W�K��2�eYSǈ0�+u��r� �����T�锁Տ����Yk㫵7�܊y!jY��݄8��NF᷒b��pB��ƪ�l���W�*��3d�\�e5h�}I��X�p?=�&!� �B\e�p*?���8�Fsx���xܱvh���u\�@�n[�j~���:a�z1R���sA����,KOp?JK�
�q�����;�9��=|&#�d�м�/iSZ�����+���f'�^�<��$96��������j��Gz��%�:W�I�z}r���������HL��T���7Y$�u�ZPlgO�P�E�;5i:��Ŵ�Q6��qf�!�l��Z�r[�Tn�Q�	.��w�`e�~~^���8������09%���O�{���������:��=�ʖ�/��e����à�n����xXċoV�hJŠH(�.�D�9�&1|�<r'�y��{)g0Q��M&>�Kv����fs�����wWSp��UH�K{x��(�g�e�"�����B�RS�`!S�M���O˵����e�|�v�t�E�g��sr���d ����Z��|J�~��;�'�˃��5/�"n�7��+t����N���7��zޏ�aGD̜�u����ƾ^.
4��P������L��ʖ*�+zY�����=B�/�L+����"E��h��o9h����鉀U��J�:����ݭ���"����37�G�������1�L֩:r�@#�6V=ϗ�M(*��NS�G��"uU_i������Dg5��y�3�y��9�B�Wyu9�؍��m���=�I����1u��?
�r�3��(C<�%dDt�e��H-!�s��Z�z�Q�N%q�E)Z¶QӼ�v'�֊WJ�O�Y��Ň���v��zZ�2Ӧ��B��B���O;_.��8����^�Db��Bus�S���& 3�+1V��׾I��`������b��AD�\�H5����3K�M�Wv�CVf����)=_}���;0�@m&�Z�t��m�S����\�N�i"+�8�o� A���q��j�W���w��t�f�N|;����
�W����@��UA,�&t����	3ۀ4&ǯ�$������fÝ��ۑA ��;3��R�.�3�8���ND�>�f֬�IM����Śy�$���8�R�"(���L���K\%��i������3�����~��.;��R�wKV����32��ͺa��$�fc�<V=ԅ�޶�?�fb9L�`�D�Y6!Aں��+�����Tla>T�z��`��4���͋�^a%9�\N�"���jt�Q�y�^�WY����1�g ��?U��6��(F����ף���@Tg;�k��\JA$��A�g�	���!<l��ŏ����$����?\��WJ�|=簄T��W�_I�����̭o��3�9�?ǢL�'O���Ts� U1�>g�+4v�K�� R�&FEhަ��GxB�s�\���0�Y;�ʋ���>6�p��6i@��z#�Qp��$U�TS�	ڂ��7>��Is�y�i��=�?����*�>d벶_^��glV�ؾU.'���g#�H�ʻ�,4�ј���� �}ѥ����G�姳�)M�qlX�t��ѭdz��p�.)�鐡�C�L[�	J{#�{�$_40�[|1jM|�|�|·�9�M0�{klݴ̇��c�%��YLS|�Y�_.�n���'��2�
�Q�J�0��?�`ߕ+�H�S8�u��T�K?�zpn��,?س�����ʞ����G��1��wˇ?��$$�v|���㻠:U��D�-#3S
<�it��Tpۏ��sI��b�?.��������]���P��nQ��7���*[l��cX�G�~'��s1٭�i�����h�w�k-'bM�a��q
�%8G3�B��2/we��Ok�
�4fc�E�_rG�*~Y9�6ѻ���9����",NPY�>��K�#�q� S�_�3�"���A�s��Xs��G�qN���������++/;��9�C"��zs�!
��'���N&IR�ߘg �i��av��<ɝ�~~H� ��*��sE�)�P.�˝8�HX���T���x��+���^���h�΅D`��� �;��κR/���YLV�M�͏xs쑀�|�ٽ솓����z~i�nX�^m��J��}��6�C(} }fmXĕ
�rs�ۏ8�i�Ub�oZ��D�@Dʓե�**DS�s�'5�C�&�;���Eg�f���l�ߊ��$!�X�M�_Π`rf���]��e�k�S�+u|����*�;��"���b`[���)E~wyS��^W���A��l�Q��n���oc��4�M�{������Uy9Z{gﴔ�����%\h���s�����o��4t���ǫ�9����c���:�i+7�����āFH�J�1�THh�ʏ<� ����4����n|���PJ��|b�5����s)n��3$�v	d��J	��g�[S҆�*���~��įކ��%>&_0�V���x�i�^�3(���U������q�s�m`Qٹ��r�oN��Fu����=Sl�4��_!���+�n34u쯔�|]@�B���P<Y��S+as�ӻ~MT��1.�3;RM�d��Z�*��� ��.6��p��/9����5��4it`>/�J��U�I�NO*}*z�)�bI.$�lȾJ~��
ФF>���!��$_���׾���΄�Q�N7����(-&���kB�-���ݬc�C�}�Ծ����N���:u;�7�1��vPL҃��:�Ӌ����j�v�o|����wR�$\1�����V���%�5�]n	�CK!���ݐs1	��<�lI��@�:���W���vzH�#\$���Y�,��#�F��EdH��T5�h�z�l׈��m�� Un
�Z5��G�}��@�4*>cz��$l6�tX�G�~�6m�(�A���M<�qʩ$����
�f�p��F����:�6�Z�v0�#��2�|X���M�[q��K�l��`�G��Q$lNU���陣w:Ķf{�^ee��(���Q&��A�8_�]�qw=�l�[�[k��q����u0�?A7:�B��l<z/ :|zS���L��Ә��Et6��|��`Q��?����p�5H���!�1��l�BWb4�mdp�1�$	��UY���T0�Z�{�z����f��oU�7�Ц9�c߾�:���\ث�`��p��4�R<6bv&��zI���q���w+�1���'�9b���c^���H3�ƀm���)�M�0<V�5�Ĵ����R��U�)�	�T�iM�eN��v�S(�V�_�A�A�`)��PJ_V!�ēZ��������Yz��;ёā7�a���!�Z̍�J�i7����e?��C��`��pc$���bGC��;Hm1��r��y(m�x��(�롴Bp�V��EB6�L2�jHk�eu�bև'����W���V�ƃ������ޢG���.��I5����sŧ�vc�C���I�3�N',�����[�e�`g������Ne�q�䍜�Y�=F_O�mŰ�'!P����c%S�8�+���!��@0Z>�:_jV�=<�r��W�t���V��d��$�o���ogYNZ��_�6K��C
���)��ኯ]�+�Uyd���j:4)ig� 8ݕ4���/��[��[�<I��-A�#����u�|~��Ԑ��9����r0|t$�-���q��_��5'�����t���^�g�Gyx�]ߗ�,��_f-T�����v`}�S�k��$�%���k!ڨkK_A3Z��Ŭ�&>(�M��t~�嫦i��l�"S`"8}$IQp�n��J8R���5�#O��m�Q�j�\|�"vT�)~x��_�����ԧw���ˬ�:�IR� �~u"f��YF��U~���[;Lq���Ȣ�p���	l	�������{���^u��b�N�}6ݩ����e�'��R�{ݣ�8�N{�$<�Ck��ľ�A�@h1Dm�F��vJ���(�FK���u�\��;my��oh�~4�	�C��*�����>�w�xg��B�M�	�Z��W����}�mק~Y}	*���5y��A�m)�o���F����!����ư7�&��7)�}<���F��Md۔1%�`�t�3���kz�A��_����U���=��&����N��z]*��%2J��Q+n��#-����B"<w?��!��F���m����7�J���%5��b;���D>�O%~�!�#6(�N�a��^�:�s�%b[���㫞O��'��yħ�YE��g�����'��3%&�KaZ��D�:;���̦�9.eE��1��/�)X�-�pvA���=^�Zi��5Ɨ+h%�;}��y��Z�ܿ���[���e"���Oŗ���l6B/�����8���6��#��!n���|�)�4ˋ+����s��J�I'�tf	���ʦ�x� �˪��N�E��BT��(gtS��%JD��z�� ��;�ȨѰ|�B6joq�"����@�5=�8ʥh�JЂ��8�8�I��I%�e�j��p��o�YK��CE��੆�R�������M7��=�r����"��Z��
����P\����<?r�j�(������<,��*i���456��m��Nł�M?����������:�j������(Ş�6���)���`$(��]We^ɰia���T�ц���%K�����|�;��c@�VmI�4����B#�YT*9.u��_Ev��q:ЪK����$������ǜɼ���4n*�	�<S�SV�O���?C;��_Pݼ���
���:�z��ph��#�<���5�ų�^���փ{̼_lF�_�������z�S�eѷ2�ȇ܈/��AAWW�Q���������<�j��k���{�������߸���`�oRt�A��td=e"���S�})FFtL�M�C��'�h.B��qS)�4*�k��cI�@TY�C��f����.WXt���U\��L�5;M��y  xq}F'U`ާ`S�H�C�G�kp�9Þ�2& ?1�/c��K^Y�[��j���@$�"_�I�W�ŝDxb���I�+�l���d����ﻠBe��m��(':��50��4y�t�Tl�Oٳ�v(��]��{ u]����d���W"��L���Y~�T������N�� .��w�H@$:ќ���}'�]<��,��>������^�Z�C���=�Dӈ7�6��a <,4:_�s͍D��Z��+0������p� 70��0T�o����YJO ��2O�t�~b�y֪����������_6�WU�(����FL!$�S��f��g
��'����j�O�K*~86���V�P�lt�SI�/sP��,B��2�)+s����؂*�%O��Y�q��ǃ��a�A!F�[�O���Y� �*3>���L��}�U�^㌻����?�^��)�_	D�]*M���a�8em�}��`n|�Hs^�N��Zm ��������Eu���5J⫏H��TXJf��'�8�;	M��o�N��Zv�y�W�dt)a��������l�_�R#��ly4�w8��Oss]��۔����8����}x��\I\�w{y0�W�"3R�{*�7+��	1�ɑ�Ws�\h�(qO�h�������m*��!`��&�����\q����Z�_�(��C%L�<C�@z
�/xխdRA�w�Y�b=�.���fu=���O�12�?������C�E��.c;�5��WnF K�nU��	��!.�}w<7 ���r�d^�1�~�d�hb��*�5㱟Cؽh(LZ`�-��?�S ���r�╠P�����QnВj�Z���=rE�բ[��:7
�)[c��&O�ާ�.��u���BF��p���}f��W��Ǭ/�I~�������',��qJ�Ҟ��6|�*v�m̲��y� y���ܳ�f���H*��
����~���0$Пy[��6htA��h���ah��R�������z*���A�����I��n��ъ.r����/B����ndR�塅%�+/`:��A�i�@Շ�j��4o�����X�A=�0��AI�[��q�d	��6H����nV��ɓ���ʰ������bvhf��������]P�*�B�UǵB?p����
鍜��:D��M�BEK�yv�N�)��.�+Ѷ,,5� dGe��q�1��]�����6b�B��u(J���K���p�p�R�-�$�+Z�s�Ⴠ%���<��{d%���-������D����uVr�'�V�^��o�|u,!��Cr4��@�<dZ��'����{�j�"��t�	i\�ݳ�T��� �z��;��Qy�[�Z���[�߫�.��"���?���ߵ֕� YX�P \h��������+y��{��5���*Pɇ��OJ�RY�:��z�_w���+y��:A	V����`�cBC�r�B�7C�Н<%���U9��c�>:-�n�+�4:p�tqf�c�ί�*��`6�>AB���f��k��m
�����\���{��W��~�fT�� �d����Fc|��Y|�0���S��Ѐ�ҫH�gy"UȅdABȀ�h����%��T8����O�ņ	��C�;�]	1A���%��RI���4h���6��i�>�\�/fժ���Ɇ�q;l������q��B�mC�P����X	�(���?��kK$�� �D���i	yb��+}��x�^SSgc�#�ށ�X)5��jFnJo������]�˺���V�t[<]0�K��k�0�Cqx�Q�������������!�W��ϫG<��;5@�ݠ<�L:  Ra���p�m�W�����gm�GÅtL���w�ڻ����� ��d#S��˜�c?��V��i}˔�dK6�/0�N����H���n�*�q�^e�!@���ȼ�2<d�\&|D�*� ��R|kλ�Z>�
�ս�\�LL+�Қ;l(m5��;"�T�\ŷpu#z�ژ@`�a�(�{���<��<�`��0a62�V��m�c6�o΂B�P�D�מí̲-UIh��~�)W۪C�߹C�5XS3�Y�����,	��Ki���Wɷ��"�Ӳ���sX��n�@��/PN��O�-���)ڼ�aW��ovr����Z��9���e��ˣ��P�pPE���4%˓X����؛�������K����ā�V�l�;�_�P��m��]��[�\ǵh�p
l��\�0�ng�VT|�̌�~�9
!Z'I�0�<���r�1B"����O�`WP$ǡܕ��-|�m��x��S5J�##�]����A<�'��pe�C(�㊌g��eu���0rʶ��˹+�r�4�A����
��`l�L���f�y�\��<�`T�l;'9���E����P��\XF�i�$B��%���y�ʥ���[�0���H}�mݞ�@:�nݒ1!|
tO;"�w'*rjE��%�����/�ӶG��"� �n�����Ď��"��8���-(3� �c�R����
����ab֚� �����w�����bu5�ŀE�P6n%�c$�S,���쎦r�[���;y��+�rN��,�<�w���"ڈ̉�y��;*Ih�H�_,���yVټi��!Q!����	��֧g�!�A�}�P���e�?Y��K��Dڙg�j,_y��8�_�����Q#h��k�G��뗪ڕόi�v�e���;�NA?�d�M�+L۾N�v� ������t�[��[N@^���'��z#��q��)�]z:6s �Du�,Nz��y ��i0M�ꃠ>�t�|w�I����\�Y����YG�q��B**�V�p�'x+��wk�1\�Ltu��ˇ��j�b��@��(x��}rt�|��̓8��y\O��"=~Qh�u���\D*�8���=�U���3�ŹR�\��b՟�-��\��������.آ��8Ǔ��YX��S;E�����e}�*kr�YJ<������j�,�������sB��Q#y���+�$��e
x�*>�]��J��t���S[�Nc������:=J�
��;젆y!R���EB�q�ץG�ʉUd�!��� yG�M��Ć�_R�հ5R���������0r����&5��;|��GmR������vW�0�N�Ӊ!X�:,Qj�h9M�F���%hO����?}�q��]����`��U���-SZ�������R��4�6�����G�%���e;D��0��$]�Z�q�{>Ň#սp;ҏ����
��U�,��nD/ʿ.A�"#�[0P��"��U$�n��RۚoM���dH���ڭ�i���k�\�v�`b'>���RTB$܌�<q��J�V�ޏ�
����4Z��Z�Ҳ��Q��D@)g��|��7�:k��	kƉ�1?��@ǖY��)�������)D�9�5�f�<wJ�6VV�����?�8i����G�F]���ūg�5��J�pjk���7L�o�/��4�M�hP��&��V��N#~-�gܣX���־�����19�=j�^[ckړ+�Su�s���_�8Z��AY�u�Z]� QH4(T�%u֧C�*���$�{�駇8
���x��"���>ݤMm�c;-�mx�~0�5,�-`Y��O�=B�a�Uy��/N3i�̄�1Ɍ�e9��P�oo���y'�C���E�M��U��B�ﶗ�Ivڹ��Cwǌ�6,"C�**��v��6�`�[���)<%��ZY*ݗg��t,'s�ˋI�:�,��Ѵ<�A�,g����f(���zT"�ؓ��k=�T����~IT{%2��v�;�Mya�U�+g5��ʐ�ӬPɝ�q��-�!����0F?�7����}W�iN<iJs�Q���Z�~�0�?�Z�pqH���O���|�L|,�5T��\���jH= M�p�T���a)9�	���:������'�$-�X`ɿ����/v��w���r�M!�:[d ������k��`�}ڛSX�XN1uT!N�iD(��; ��B8a�#��3'#)���
�Hcж;:�=W�hV*�y=.���.탘�I9@Xq3�q��_Y�41�Z�ࠐ�;�p2����R�X��Z��S]��^�G����,x����d;��%:��M��prs�E@7YF��T����W��j���o��a�9�j����Ǌ�ٯ���7 +Β���8:���YFq��ʡ�b��O�B���B��S�4m�F�S
��ŭ�1=�<[�C��W�(�WJ��O1[YN�J�%��jl]:S����>.dc�t	B�tz�]�L����p��e�tn�B[p������$)]ƄC���?��1S���Fܞp+�H��Y����o�=:�.��O/�@�S���'fa�"[�h��~Ȃ��m|� ]���=�zGw>ɡ�N�r����bEN�w���җ��ؙ�T�� �ؾ�	���eD'h����I����-��9�u[d�
����L��J�TV1���z����{��� ��=mI��Фm��@�m�'��;��>@X��_e%��������l��o���+���ny �����5�E6!$�_��,H���A�y<���ϝ���K1��ն3����_����k&�q�疈��g"�Ք�)�RR��$��Br��:y��΢9�^,|� ���w��#����m����_h=���A�x�M��a1�:f@A���& #,����{��%��8��qE����!�r�i1�S�2�E�
e��W{W|��t\�X*5 �(����8�Z�2r�7˷}�\S�y�R�P�FU�࠾,+�FG7$P���������,ն�W���۷�{<�t�2�9+�>�����jui5}�~$=�X��(��Ɯ�O``���	�c����@�?��������=3��۹i�.ǝ�����=���w���5.����ߨ1��
����h�W���iag{&4m�
�7�2��2��R�\{���^���HDs��(�w��`�rS��ҍ���1�(Ǧţu��/G)�܍]1�2>\ܭ8_m����K��p�I�f�˻���Ő��ƺ��1'�;�6S�_L�����B)͆S#_	�.�M�h���<Ȱ1�[!�q��!C�a���ȱ�!d�8F/�����`3U1����uH~{�I�6ᠡ��R,c������#��|h�:��W}�����]Ru��:�ee�x����ۭ
<-u���+�X�(�/�B:����_�l����o�nSv����;���Aq��,�a���o��M5#��@�[xT�e�MՔS�����W�n��W�ʳ>���4i�}��>�ӎ~�J{|�,�:����^u��i��*J�ì�@��s�tK�8Ou\8�e�Rr_�q.��y�F��⚏�3J\h�����D-�a�i
{�P�+���}�8:��h��@3���׿z��h�֣���k�h�ՂM4���m��Nbl��X�<e��$���ע�D3���������r�����4���`zt�:!@�>��?�WQd=xA<���Aй���i���Ӧ�s:I���N=Y��m��a�(�y�9D'�����k&�K]��*��ȃ�֟y(��c���w�-��$�b���塻�;"G��r9�Ԃa�ױ�av�;~}m�VN%I&-���� t� ��)�H�-(v'o��]��&�l�}���I^`�3դ� .9�?�?��<���a4+!�OM�����}�J�+�y������k���g��xHm�"��^�r ��G~gNU�-�Ŭ8]��r��u�|7�%<b��x�� �D:]�<�9��%��@u��oc"`�aRTs�n�w={7g�`� ����x���L�������	\[�D��#�R������q� <S�,^���N�	1�H��++��X�yzL�� 'M�M놺>����G���*�� C�i�s0�i����g�[�iQ�19�k��D�_�}�E`Ky��l� �Tf�@���4B:*e����\B��aȄ��'r��$�0L�V'3N�o���=�G��L��ݐ^��ۆ��aٲu/�X���d��۔�AL�zú�,���!M�#�^��U�����:�ڄ�Pц���� ����p� /�{-�X�DL��xv��hK����;�t�ar��3�\�l���j�b���/�[��BB�xi�SJ:�(���^��O0n��|��,��h�|R���:�����,����5R̋���G��ģ�����*��i048�I/��/m�R߂f���L�"�����`��\?�p�C������\ ���M�Q���

��q�!d7hwoP#Fx6�����ʔ�P2۲�}����i�-����h����"hvg��,٘S�m���7�ʼ�D�g�*$�08�.vO5��DQ�kM${1���4�l��d�ZzC"�O)N�7k��g��{���=~��Ck����ޱܗ�Ӻx�:�\eb�A
_��</@7W9y�9�G-c�� ,��_�̳-���	e+��%Ú"&��W:�#|��)K��	T}"�|x��R*	K��^;��,��&������1Xie5*��h��ۦC���7�� 3"�Q�f�{��G��)�7��)��eĩД��0N<w%d:I� l�wT�=���4������A,��.�	;a偛�?a�zU��]�3F�]���=c�3Ֆ�`���Ԝ�WJ�����A�c�")��B�{���"!b�������q�%b$	d#H+w�F$��5����HÅ��wj,��w �.V-P��~�G���\l�	d�Se����UA��R�Q�XyG�r@�}�O�~?�'7��-(x���O5��C�=@DC�_�pCBFw�R��;�ٳj�����oH�9�> *2�s*�\�,!�Q��OQ8���{?�=]m��4��i��n�{�&3o����L;J3Ǎ<��*�����6|W]�F)�4��$S�&B�l��#oF��f[՘֯)X�j�@�|c���z��5��0X7C�Dy��j�j����#��S���h�w/�V�0�T-a�ZU%C���iA���������8���6�5z���Whfš�l�]̐�I�0��̰��;	蘃- c1��5	C�U,AWp=@������.a4^HdD�0L��n4)�u���s�����,3�o[�	Ʉ��bLq�J�4W��9�<ﴐ�( r�$�|;d�D�����|%>�����vK�c����C�wy��
R����f7c1U\���	�V\G�>�0�ʋ��W>6W~=�:}���gf�I�蔉�AT@fӒ��˪O�{�ÅC���l""[��y���ɧ��m��p5�8LM��;t�6��'�\�������jT��5a!x�~`�d�����4R=�^o���H��� &��$������Yo������׬\;��*�q��ve����)�c�6�	�����,����=T2&���t~�������Uy�j;ӤaVΊ���
3`su��C��+�ǧ| ��7�A���L.M��b��s2#m�3)1Z
F�.B�����EZ���0u��\4�I���G?�ub�����j蟓�,��x�0��6E�^�� �����4�a�$y�,�͸<:�uS��:O�ڦ�	��Wеhb9�P���:p�s =P?]�q�9��S��6(�N�+<�'��s��u$�����uh^h����#p$�<��>�|\;���T��y�&	��n����4w�V���F���z�'��+�WԺ�H�}��˦���;��i7|�g���)�ź�OjV"_*-m�u�^���18µ�w�r�}�� }T���[uA���בҕ��_�G!7�g��;�|�Ti'����x�����=���z|7�8g��,�y"���r���_��ថe��奋���ߒ,d8/�Z�#�Grߜy��Gt)2_�?A�\�Xۡ{j��Q�I�`�p�Du�N_�C\�5�5&vB&�����U��?3=T�B�0�C��&��q���e���47sP \��:�M���h(ꌃ,��i�7;e�س���X��-�hb����S�&���O�R�+�k,Ǆد`�8�K��kL"����{����Ƽ�X��͟��?m%�Lx�n�|�)%�tӰ�g�1>@�N�=w�d�sΟH�d%����+�F:��M�B��Ȍ�P�p� ���%��	ۏ�S�ڭk;�<���8�*г3&�/�-B�|(Б��N����_�k�h~.Ά�:�
zK��g���z��U�fqRⲊ�i�q�Jl r���[EJM��[A�ؼK��c��L�W+��؃&rP�d����T���w�Ƽ���9a�J R^
��e+ؖ=� ���+�緟'7r�*���s쌿0�M�Wq��i�f��u��;��}�,����R��PC�$��mSc�,�����EQTmfU�د���J�߁�C��M�M�)�n{9���>�ir�+��j��W�dc��������0
�1���vx/����� ����<��]�9��xu��#D����!�E�G����]���y���yh�"�⟆�5/(]ԻR���̋؛e	�V�6[,a Vm�J]_MA��r��|�����Jq�$8���X��ʽ�<0����?�`���r^=���R�n����h�T���ASt����_��zjD�M�y��bR�Y�r���M����&Ϲ�fʵ��\�8=k��K�Ỗ����y�_�LJ�
O�Qrm��_Ff=�X���l�-�:�o�ПM���O�ڝ& �&S���\�9��n���z����jz-,1_��G�%@d������ ���J�������^�1�p*� 1�6mĀ9I;�Bm�����4OX��EG��q� ���m%BXo�ly��4�8�(�&V�늘���|�ey).�w6�yJ����}lmahiڋr I���"5�#�	�q�V��S�&��	�"��-~5/7"�y�3��Y�B)@�t�8q'o��z~����\���hurߴ'4���4��0~'�j��I��xmq
<�`�K!2C�(ﮒ��eQ�8.Nά}ߒ��9R�����7PcEn���u̜0���<��	mv`�G�6���������J��͡�d�H�XҘ\Y�Ў�H܃s�%�,BS�j�W��a��5X�񥘭
(�f��߽���=��� �J��d)�Zi	�Ĵbu��,-�����`���D~�}�j�P2��Of���mVo�a-/:YÒ�T�U����0������^�H�rQc��li�%Yv�����9Vy�x�3f��^\T��O���N��]S�����_r�ͤ�"K�;Kw����Z�4�_��������}+��`	��ҀJX�_/�q�d����	E{�G$kjʷ�]�F/�'�VW�x��~+�]Xe�=����0JGx*Gݾ�l��"D��}���M1�a/D`�Jh��>6�U`��E)�Ͼ�����E�=J��	�LOV���O)�8M9���~�Yε�ZnE�]�u���/�:N��F�m;�^�#��l����c�*v"�0���$��d��9'����lC�Z��e���keD���s]��~�}�I�o�
�GO����ٿ��G�f��򎥪8n!\�����gP+�$�A$����%�K��o�>�qS^y:����1�':�k�%�i) B�mNw�s꧎_�z?szzNjh�a�[���WA%r�ٯ�����	��.�D?��4�B�e�b�dhm��':+Ĕ[��O m�R�7��BL���`�{}��l�	��ˮ��5���&�"WiԈ�}'�g��t��[ul>���N����G�m�A���s3��U��7��\�'�����~k�9pvuRWx��/� ��I�?"1�%��gz�=���52�.��C�=KIT��|�?2��Qy%R��:�7/���#<��j���X+�=��J]��wT@��*w��]^�����Q2G���{+r�h���j��E5g�	��:�*X$�,ɕő��w��D�%�ɇ	�׈TP<�iU4Գ@��*�k$n��%(wd��d�Fa��������VF�;n]��2S]�`%sC_����w�َ}A���`�R�����m�����:���!'����AN,�Ee�ح�-"в�=�9Q,ơ���\�_ё�6�����������Zy׾��\���J��.h�˭��	����v�S���4��٤^p���w�����YS|�3�D�E��ɬ����ip@�l*)���F���Fl~IH�M�I �v:��H�S�X{��{��a��u�[��:; ;UdA|����H��
:�|Iq���1�>��(Oz�sP�ڵmQ�$�A��ע=E!�z'����Ќ�1Jas�D� �٨��h�f��=L����0ןiE��fƬ!P<]�AY�"�i��#�A��.|6�$"5�]5�:�i�/lI☸�h/�cf�?7��r�U|�hP��s���b�|�$�
i�FF��N��O�wƖ�v�Ҥ�|-~�4�_43=�U����n[j�͉��2�o������9J[��ĺ �%�/E��������+>���%��=W~�6ٚg�xAr�нE�^Y���LC�!�D&�R��1�D��
�g �j���V��^.�J�e~]�$)N����k���`�1�=�9����a����i�V�n:�1V���Q<���\�,]�Ѕ����R���+�*66�p���H+�������[��WM_YӰ��l�hԎ�&���wr���O~�;�T�}�R���g���qK_��6U*;�N����KYr=��6w��Rl�0ۡ����NA��ԮB�%�T���_�`�-�f8^!��� ��y�;|���������X�Z�$w+�p~�P�t�i���-�r�,�ˉ�
�3VO�� \��B������V3�}��e���u�3&�l	�ޖ��]���#�;��o1��k�{l[��U9��/��;��Jڠ'諾��7S=��c1����L֘=3񭢲�hg�-��w[�����k��4w��>y�U��4pS�-+r��<�?Si�1*�b9�8Zt�@�x_ͭ�Š�'�n��eR'���?�P�I_�O���-A�	�WR��
(3]���;�?��u��	1��%*��Ő�~#���I�%?��2�m�G�ޚI�T1^̕�Ф+��hd���G�π�i�`�U~������|��N���]I�C��ۉ��+b&���@�A'��`#5:NK���X3z'��u�M�^��K[�+r�Ş�5Bp�bǘ�W��:�SKB�;�/:0�����1�igp#�0��x�]����2_+�^S���P.DN�>�MY�_�sF���B��<ckҀ�V�}��)�SSC]R�$��Lr�q�*4��d�Fm+E͓�^@����VrUE|^���`,�&�H���̰���}��4.-HWQ�É:Qn�o��^�����;D�NI!���$9��c�ű1�H��/쌏�����	���� ��T�&`�l� ֒���Y�`�$����<�����:0�Ԉ�w�����[�z_��{ �0�Z���	M�,"z�\H����D�W8x�gf��^q�&T1
������,�Mü�ҫ�`.�YK�$��Y�'a���/J�n��] ���Q�(@����v^�K���쪾I�}Npj�K@.�5�e²�f"�5�#8^@�8����pm��a��N\2��3��l�vq��lz�g:�K�o�:5�}f%�v����h��x��!E�0���6�^@ _����R9�)�[o�z�x���U�D��n`[�����8
Mo���E���Q�J��f��|Ҋ�Ϟ��,W�7�c�q�2�L�]�_p"���� ������w��+\��rsZl��<�U��s��Ac,ͮ���+;�D��X�7�`�UY'skx�w�o'��/��'���b+���d����/C��z�B"I��6/��4�
ԑ��L��Yͩ��*�G8
�0hJU�=���ɵ�I�O�>"�P��Y���uM��Ne3\����Om ,d�ƽGr�(B�L]Y�Ȱ��Ps��,Iub�x��RA��B�
�cnʈR�O��V�����X�p��ڬ	U�xX�c�4���*u0�d��m/$�Er�e�:9V��G���͒B��%��F@`e[�Ӆv��x���YM�==^?U�6���t%����G�y�9�;��i�[S2�l�Ԥa&���TN��}�f�:`�J���^�?���n=Y~^@^����U;a�I��2rw��1��
��ۭp����k'��zH��hZ�z)Va$��D�QK���jS��v�Q�L,�?޿��w��͑����/~L���~��� M!��a�?��.��{8�7��=��O q@H~��԰��#�`���R�t�����F��aÈ�c�'j;R�+�L]���ȇ�ʮ�RҮ�p�hw����)�S�=�U:�Yt�m!zVQ��^?uϞ���ȈY1F��2���c�_���?�dd�� �8�J���h8�{�27<�E&~��%�K�{Tr}���������}�9�k����.@�6Q6�N�TD��/�<h�j�WU ���c^Q"�R�w�����\��e��I31�Sm$�t!��b�Zh�x�۱ӥ1���VӂD~&��-�`Iz��Ȗ��M��y��%[/��Bc�}���
�Ķ_��Z��"�Ɣ{i�ǌ�a�?�g�(u@�+����=�V	g,����t�:q��
l&	s�q��_{�!�ZhY>qӂ����t�]�7�]�?pEMR�
f�!qvIyN���k�q~&oa�6MأL�0J�\O�����M)	#�����ے�Sn�qJG|���;\�m����}Zvc��v剌y~n@�h�ӛ�?�D���)%#���V�o�<R��&[5�@��4���ۛ#���)�ʴt	=�m���fx)����������i�]:M!�a�%䞷��l'1���>PY��.G�fO�/��3BGD?�e��"�ɳ�[��+#��퐁"�x���e�%3��q��v���HD%�Cy�^؊��Eib��-y���J'n�����0g�RA&�8|�ٖz>h��i���5�]g���L#�F�Ǳz�E*%3C�bj ��N�u�O��k��F"þ�O�vs?.C�k0���P�b�L$&�h!x�l���wL�
��l������-e;m�/���Ee���6���~㳾��;��,�3�W+:�޶��.�
Poп����@�ޅ5���5�11�߉����m�F��yr?�<�K_z��g�kd��ζ	$619e��� ��$���m�#��>��"l� N�aa�=,p0��8�$�/ u�аA\l���̛${��F�e��g=u���@I���5�ViL���z{�A'jBj�����ط�lM$����LK8�\?�7���u%V��0��CK|H��-���|�:i��B�G�?v�B%��6�+|���f "�}PW��;�(F���8udd�7M�Iք���u��2�pv�x�H�z�o	;�϶ڨ�&�|X_���O|b��SIvE��ѽO�h����_gQ��}���>����Wcs~q�3���[YA@���m��N�����AM���^�D�~���w͈2��+e���Ne\�zm�Ф�
�d�Ć"��$7K��)�_2ٻ=�⺼G�����$���4z�����xb�]s�@�2����$n��9�*)J�L|���9� �-�Zk*��E2����*�M�r*k�������Ηu�{ ��XI�iI����Lb� ��E���Lx�絈CzAւW���gc�+!������)l�����w���rt����K ����G��ZOo����_:�ظ�q�4����0k�wd����	�g��� ֶ ZX/�iqi�Mt�V�V�]F3�C����hߞP�!�Pr��7u�F�t�=�m�~�a�L�c�|�蟞���.��}�>��Q1��Y�D��lZ���#�H��G\�4�& wce�9a��K(��B>�hDFm>mE��^7�Cz��1�.Ӷ�S�G��}2���*�T��� �j�Ķޫ��ZΒj_�=���lEY�rR�^R]�X�ۖT������/\+4	��}�e���1l�'�ʝ#RɄ��������$/�1T��v�t,��Ӹ^��rd9����T%��=h9'����f�n�k?ˇ2[��r���Ѡ�L:�XL��\y.hL�Ob�_�˽�Z�۽I��k3³a�.�W#	�"׽l���iAL��0�נ��~�
����F��+뫼Þ�����j���b�k�����$d�_�����(ZMٶ�Z��u{�6�}.c�Dro��s����g��I�I�T�XY���Г�ÿ�N�!w��	rXu���2g�/1?d/��c{;M����>K��Qo'dԽ�j
�K��$�Ǌ �B�A��CC���Ǭp�W���sc��M:��^����"Sw�4%�N��-EE��Ԗ8�9n����^���H8�ׁ�WH+U�^�|����S{=��k?ǭov��d�)���2��嬑�2QFzk����JNL�uY9q�6�TlP��~Y{�g���Q#]ܞ�<�^�?L�|$?k�m�[��hʉ���H#��y]K�3N-����T+��٨@���A]h��T���gW����q#0�`]Z��Tԍ�.#4�.���>�V��$�A�iM�I�Hb��Io��G:�T��u���1Iܹf��.&pr-Ǥ$3��Cs���>H@��_�a��".�,��͋�O.���o�1ɈԴ?���U�G�;�E��
�KO�zψ��`T��)7^͋'K�$?W�:�do�_%�|:E���6n�^>�����Q��6W���0�C�w(]Q�׽k��� ?H5� �қ�W���i���A�w=/�~���zыq����=d-�h������*g�uQ�0r�pB�s�xJ�4����g�
���=V�3nl�*�ӄ{�A����kׇL(;y0��",��T�<2��%k����EI��0���'_�z��*��kO�V��K�7��Y�[T3�����q�y�z��U�3��.5�x �ސ��q-�O!���L���`�d��x�K0�ӵ��4E�{3��/��c(����r�A���S$�B��NvyC9&�D�ջ�m��-VˀI�N֥��pLI��1���%�B�N@�fq[��1���mA�\^/���rKR���Bå�Q)�~Md�>�Cw�F<��)&�:,�v����.��$s��FK	���5_�BY��\�S�W�5(�7�M�X�`�>��w��F�c�����(/#�ux����{@HM���i���V���TV����a�Nvv���%��`��� z��� ��Q���ӓ_!�K�Ü0+c�1������s�zMm���F;�����O;VX�@�I b�ɖ���P1�yFN�$�;#��5�4�-�A���)��y���V�;Mܣ�3R�4P��˧��f�-����uw7|a�yp���?l���<�diu�A��&ȇr���  �#Q�[���Pg����.=m��9*W�7LY[tM�N�AD3�|�Z�{x�G"~���X8\���P��l���W��>ւ���vC�t��8b��{!xH�*oߌ��
�[�r���nw�̶|u#j�8 �[�[�ۏhO �(`f�;��$X�Im��Z8��e25<�:��������H8�E:1�wd���(�+�+�=�&��q��<�N+�NE������a>�4�`Zjӎ�z�cϓ�m�@eI�wcq�� �+#����brCC%:`�I���7I�B�#=쉯/�I�=�*l{���Z<���	[5뙻o�`!vͶuN!�
��a�'ՊE'޳����*1ͺNNF��MVf�tۍ���4����W���FS���8���DB�rG,w�:�e�@�"m����D���L��(�W��r骟�Z�x�ţ{Υ�%�Ov�������-���@����M�2�c���A,�����1��a#�.	��d�f?p�.�M�����u0G%�z-�[;-@�͈+�E޵���[�%�^�A�
_F��iF/�=${E�kn�8i�����_�'��� ��ڙ/�lU��~@�ޛ�W	DԱ}^��x ���J���\����n���f��w4A����oC�͇�Ya��T��N��/HAO@KK������Y�V6�s���F|Ci w�~�d�H<X���4c��/S�r�cI�:����sY���]w��?��@��o�9B�e5����ٗ��aaQЂ����M�휉2Ҳ!��QMxa��/�;������*�_�F�>%y�
��h�8�:fW�{�a�T��_������D���
��*�ص]d?��N�X�u6�,@ځ���;u�~l7|���)xS������閭�=2.M;U��z�p�;�/)���`�4l�|@�]���|+i-eQ�A2�>U��])�TmD�>@��v~2С�b���g��w�{�%��Oe��^ϩP�n�����"��ub�tY��to�m��}��Ĩ\��1�ՑOb�[[̾|��q���3��?.�zr��I��hƼl��>�/1��$WU JL;mB����t3h��ޚC���]���+��:�����7�ޙ$�́+g�;*����C�S���e�p/y"�S1M-��<��z��{��[�s|��2��c�'+�\{{vr�q�f�6��e��p���,�y%?����� 	׫�縈�*�jL����5�HЬ;�K���Jy�9�\�R.��Nm��̻��7L�b�-dO�� C�+�.�yL.baoL��0����rS�/��Q��^!� ]�f�mY���ܔ4XÝ�(h?���t�0Π����Efwl��}'�w�(jn�K�������ԥ *߲ѣѱ��^��g`��I��zG�a���N��U�k�>N�0�~˃�M����/cN:�Z��k
�M����~7��BufQ�K�B)��T�o��JwS���?�;�[�V�\��9�a�g�%���C +y�-`�l���3�`�O>?��Uk��`ȴ�w�D?�I���U���R������D�9T�v+W&�A�����Z�t,h`RP�'#�{����,�uțɥ2�L���� ���m#��Y.�K��)�� �X*z(��^i�â�7T��Zh�q�q)|܂�3(�wܡ��%�r��w�b��)�7��|K��;�Ke�DrK3�V�P����_~�&��4疽B�*s�J��|N
A54�M�(�����T%]EэP�X�>��)��*�َ;~oz�>�\G/�5��[�wy��I��@��1I��H?�^��u��3����Xi���R5���mb�w�R��{U�/����	s��Tcz�^q_>,޶I;q<~�n&i����0�\h�)o�'0{�D-H�f��3`�w��8�� ��>X{�,_���y��֩ 냵)�+�9
�Nc2�1ޞ�A��}��Jϻ���f��jٿF����#�	I��J.��u,t� W%�ADR:)h�6a�!\#'^����G�<	�A�.jz�G��%�j.E(:��r���0m��@�x>Ͻ)D5�����~��S��]��$��/��C𓁲:�nZxC�"x~}�H���<V�MAb���˦(�֠�ԟ�G�b8s[Ai��-���J�3��������٘zǬEH�e):=��
�?���V�����J���tΩ$�7x��5OG8�B��N 8WVs�[�"���)��&ग़�C:�E����~;5�H�uX(~VѴ��}Ӏf��W;����ee��х;�R+4�ø+Ҋ ҙ��xg9�.�\��>^2֦Z'��ݔ�6e�a먙7�5A�������1���i�+9K������%}�P�vC�����nt�Hy�]H®��g"I&�D��9���B)u����AX(h���T�bg��"[V뒢�:@vqw�L�T5�bX	��I<>`>H9B�N!���-��|]c��oٵs���h����sj?7��/�*�D�&Qr�iVW���<�/���]֓��dql�F��é!� b�JKr\��#w]eV~`�F8���12t�D��a�ƖdJ�:Ek� b��N�6=,�	�R���Kq85�ˎ]�������>^-���J�֋�o�p �g��6QW�p���ϰ�q'J�r���%�WY:͹A�}Qv֊���v��=ũ`�g�!����Q~�bZ��,%6�1:��ܧ��5�o���9z�V�Na8�[�br�����}� N���ST��P�\�I3y�}
@�`�^�!�M�N+����X}��m�!rXL��+��ؘ.P�g]�����i=���2V�-��#�5*����++��ye�r����IN�,	�`����*��.�ͮ]O����Z3v ���|v�*��8nb����b�X\�Qn�4����WEj�m�\�}EEb�k0B� R��:�	�bLu^�9�n�!J�"�,�Ec+���ӌ._����̌p~��O?�xG���fl���߹8���d���9�5�/N>�K�gBH��Pu�1:�0�
�!��P��:&�8�TEe�Xg	쾶E�E����G�vf�ڤvFk6�R@Sی��"�úP��N�F��^y4��<n�b�`�_[D����VlzV��:�9Q!Q���0�&���T�����9�r�k8T��}�ղ���F���I����S�m
l�foP�4�X���0n!��p�	��Gm��I;5�K�Z'�G� ����\Bv_����:����/��r� P�C�;;�a'+sS�����QӪ?Ӱ�lj�	'�,i�h�['(F�m�5��{0�?�D�n�~6���o1��@�R�j�/�5��܏�;�r�)�3uƣYV��mᴧ���jXw0(�s@��E�Yւu���5@]4=�����
 Ss֘˔'5�Ha�z�K,21J��:�!�ڬ>�2o�b�Eq����\f&N5�/�:��{���޽h��$Y�nEE��� �M_���T��"�`�<�%g<L�<`U�L�솗lރ����1�]b����P� \��<��� ��"0�h:�> JŬl0�reIw�v�	��+N����}���X�}���		�M�KԜL���=w�d�f`�q�#%����4�!l�s5���|�����6�����Ms����#��R�WX�>[���S.�E|E¶.���k�q�@/�Z|�~��H�nQ����5mt/�_�Y��3�H�������)�����v�9(RZ9=�91쳐V�S�	�z��Â�7�����^��.�/9p��Lt����O�m'�.�? �f�u����uFcS��S/�kuu�<�͚+FJ���ҏ�ҁ]��R�{
_��Z���_��;�y9���s�����L۪b�3�8��6's����5�������YV��j3��ϖk ��`С���o������LG�;ك>:�GK`ߠ������;���8�u��# ���mq,����+8��xv䭹��2�H�����/��/�5����u���^��o��L� �-É՛�6+e��k��o��*��0���0Zć���Y��CnYփ�c���P��Օ9yf� �\�f]=������T� �������j\���]b>��c�W����E�d;�Q�D3�`9�U؊�+$��.�1�Z@�5M�wG��6\�]��")�p��$
=`(�6!���xL�>11(��InŤ��J���e~F	=) �xJ���0�8ho=ٮ�e˼5��e��Vv���@��X:�����,�$=j�nFސ��ϩ��w�� �qԱ��&�d{i���u�~�6�Ħ���n33�ޙl���u[_����~ ����K�|?��P�����61���>Ԙ�����/�_���$9Y� ˠ�H�m���K�q	�ж���ZҚ��F&�OWR�$o.>l���#32��)Ywp,צ��.��=�W�/�	@����5�d-t��\˓~�m����*�6�O�'K池O�|zKӶ��h'Q{y>J�.X�|�53b�)u���5��t`]Ag��U=�!1wo�~��s���z��{���Ek�}9Z�t�������*�E�yiQ���.��ˤBY�|��lЌ��>45��-�;Ɓ��0@T���d�XM�M�=Z�T@,^S����+��2m�߶��m��F|w