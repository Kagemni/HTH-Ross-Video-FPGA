��/  P"b�z��r֪��i��
��q��n-Z����Ycg�D�ڜ �"6X6X)�ϛt�k�����m�a\8N	�AnCCe�'�Վ�tuo޴:!���X��,�m��������z��c0mg��V��(&�j�dW(��յA�D#���}Q ��~���nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n�W��ߌN��5=�8�:N|���gp�P�ظ��U��)�& g�J����[��kC���RmIOʹ��Ut�~u�4�s�0}���X�5����M��Һj^����U#cۦ�2��֨�����à���2S��R�UɆ������k�]�!]?��śO���k�Q�L{4�1� (�7cI��V��@PH��$9��ֺϣ
H	����?6cI���`6Ş�U���~�Z���[��H�G���C�g'L���̟=M2z��+"B1_�ܦ�1��:)3��=�r�dk�f�жK�3j��b&��	n��2G���T��W���']2�,��]%*���T`#X-�{#�bE���1�����Q�L�-Ҙ'F7��ﾄ��}ި�X��Q�E�k�NS�r�$�t -܋�+��c�2�����řp{�
����us��u���s�B�û0��e��I_���1�x�ƞL��S��r��UnTX|e�Y��[ ������	�z�V�g�qF���L�ȦAQ�C�=��R��C������-j�'Y�s@�
.��%�k=X؂d����r�?�)M){s,Q�Ћ�Zq�{��/�\~ڟ�=�\�����(�>��C����\\�\�p iG%!�/}�8����� �<�\�ɚb�<��>XE��ՠ����ECe����vl%�x�:oױ���b��E����K���ڲ=+>��
�����͈:'�@B��o�!�Č�?�I��k8���Q��@�����3��	���^3q�]�df�h>���]j����?�1�D��b��vM�gC���Z�����R��$���~�+��T��C)1�tZ���D3�	*u�����oVG>�������3��ܫ忛T�E��)�u_i� �<��t��6�V�ෛD"��C�\�߰�g�[x�
�+�U� a�c���踾L�$"Ҟ�\�o�L	K>s�Ɋ�e@#w����A7Q]0��+q=Ⱦ[��O�l&b>�Zn�c�B�0��|nHT*�& 6e'�v=P��/�H9H�F��{�������i�W�!ֿ���v}s�����A�*lB��~�L�ӥ�z#��S�Qש5MP�0xɠ�1��u�������u;��p�D@,�qH���)��>��
~r8Wg�����yg�=ߥ�T5Q:n�fAIc�Z�P=��ͬ R�K�����'+43L�U_�]֕&3���x�f������)o�N�6M���Ab&�X4*Si�v���g>��"�|!"�W��H�d�%�M�\����l-I��h��
P{[����d��ޯ*:��n�����]�*���H7hyBۑ�R�`�g$lEt�% �V��ա��95�C`�K���L��p�5l�o���!�/1J�<��:�T�q�HDb��Aⶄ􉛩ԉw��ǽ�i�-�ĹJ.�q�K�j���Q �U���瘟)����s�O�>��������2P?��t�2�痿�����נ��(�uj����fJyV�4��	���N��y�c���p���3���ũ��Y����'��JJy�Lo��W����g�(Q��;<��q��_@'�J����[H�0�,�6h��������EF��̿"�< sL
��g���g��1&T.��:A�}]�Z�� ������K�H�N�H� y�4_��);x�g��q�'&83nG!'*E�9��҉t�tj|`�Po� ��Ȏ�|�Ĳ�W��t�������:e����m������Oy3�B�4��w_��&/���~�Xni�����ʃ�#Ŏ�I�T�˒��W�}&'�2��\�Rj�nJ(I��\�s�O���'<������6����؇��V�d}BC������� й�JIN$B�O?weo��҅���vQk���l|<jKyKC��-�bM�ʔ]��Dc���D��QO���Eˋ��Ź8��6�����/)BWj���:r�.�	�A���c%�DtFc9咊�@8�k�D?���6�5�^\�(Ao(Bc�d��KM�Ls��-Idܲ�e�;����O�cM���q%`�,@�1�� �Z�SW9!49�{�>��̒tgXY,`_N��'_�D�>�Sd&%�´�({p����D3�����:|%k8P�뫯���Ph�ɉ)�1�j~"!��}��Y�S� �d&"a
����'j*���&��k�v:	w�4:ˋTY<�Nt\1sq�X����l՝sc�#z�=��e���Ʃ�Q���tg�KF�@?p��-����}酕����YS#����1�D�����]��Ek�[K�A�A<�+�8W�����{�/����)Q܍�)�`�H���"àa��&Nߓ
����2�T�=�D(�m"���<tB�^$D�F���� ��dT� ���֧��1�@G:�3Y���STN�#����t��b�x�DTU�������7�=�p�>'��$'��N��(�'g�\��Hj�Uf�wk�_zH�]�o��7'�<Ɓ���
�z���/G�N؁NÓ����Hz�R��r:|�O��m�t��κVx��El�����69_��_�6(�[�lZ ��A�ËO�Es�S���=�D�LE)
�z1������	l�.�;t��V3��=8؅c�p��Y^p8:G���ܒ�.FY���cF:6|�7_���9:ȡtw�|���.�0^���^7����f�S�$��r��N$�3�TZDT^��m�]~��~Hb8�b*�ج9���x����P���� �ԟ4���̯�Qk���aOY�.uЦyGa� �������ҍ�K�y"�p�ߔ���/7Fn\�}l�L�g:�������"��7�g=xYq���S��&�R�D��H%�v0� �p3@$e>��nZcnd��n���|4-oak�6�2[h���F��ݝ��bA͞�f�Ҽ�Ƭ���׵7�1K-���H;�R� (���܂/ ���EȀRB�l��.�K�c���Ƌ��a9#!wQ�8�Zc2Z������Y:���b�F����8,�yU������e���ʅ��Yq��O������Æ�Y��A##�E�t��aKT����I]��˳�����d#f)��텂�/�;�i�$y��n�����:R� �C��r�^J��֯�*����\n�C����W�ixE��z����~�E�U��]5��2����v�K�/�p�R���{8( H��dڡ�ɲlﶟU�¼���ߢ���M�-`$����� ��i/x�7{A��gx��H��De�2�drT���S�\�ֹz�$�ƫȊ�=��~_ɦ�#�G6�=��8��3/�e7������$`��$!����������T���码q���:���`��6���/��U@��*~�(q��`≬�mP3WT�S�XED�&��\nJ�ȆZ<�J*Y���ٞ��h�p��e��T0N wh3�!%dYP��%�2���s��&��r�F��o78��Ozx9z�*=���e�p�Cu����`ܝk2�~�s�q"}��!��g�G�7�	���%^Dgp����Q�o�Ph�ߔEd������n!��Q	� R���و��Wz�/�j~���
�7��7��5��x����2�K��B�����%�OB �}�C ��B����p��i�m��,,����f�Y�k�^-�,�Ĥ��`]j0�(������p�<��{k�
~�,<��Q����{�����R�+��v�0l��y�{�CRI���u�mv:m���'w���6��H��Fɱ�ޏ�3�����'ǉZ,M�`d�8�f}}�������&L�4>��',�@�.K-Xu�?�T^�
�q�l����udhI����z�>���I�[Ɍ��{g0줦��}=ւS\��s�ӟIN����5|�����B���lS��q݇�N�>2.�6���#Vu�#��f2n$%�����+#�o:�ic�]l�#��[E�18�tyB�3�	������M����N��.u������d_r�N��\�b�\����)z�Ud�7C?iap�q��� �J,(^���X�!�Ao�0�ʂ<��Z����~%�qW���&�4%�A�^�i���kG�s}a:��b���ɽ����Iq�A@.�E
1u���%�.��vd-3V��:�.ڬ\D�T �ƪ�:BN�^4,o"sAaM37�-r*Kk�jln��r����
�W����A�B`�<�W��٩�6��-��b��j���I-�����yB�)<_»\q�h� �GgfQ�G'��N����wx �|Ư(s��m������f��q�V�rט��>�Q~�)���WI8aId�Jp���+#<
X�+kAI��)�M�Ц��zJ�D,M�o��*b��6i�����
�\�v�С��a6`��5a7��Q�s�ϺO�����#s��=�����[F�Y}�'��m���>߯\]����sB�{J	�����[�S���XM�6g�`�6�rٕCke?\	�*CG���N�1�,����5PN�l����nMt�����q�텁3��o ��� ��HW$��lD=zn/�m6�gQ.jG7C\y�#h(a�ߐ������=�����xYŔl���>b�����ܚ��3��<��Ïu ����@<}e���E%�z4Λ�E����,�J��38���������^�w@��A�������4l��"�|�N����hp1P�ט5.wf6����F��EĪ&�������ezl]���"���I�+#��TYcs-;�w�
���t�p!<&2?-�y�r��a��t�Jc�r���h��&64-��ڙ!VE����݄&��Ayf��pЅ%�e�� k�����rn���ܢF��P��Ul�� �5(W�&��;��h�J`�.)$&�cq?�)�.��)yq��l���w��.�I޵�L�����@��:�O�4nΫ�(�`�Gp6��4��\��9�`jy��#�y=z���h&��b��.]IV��eԚ?܉���ưo�n�����Dԭ�ā����v�z'��H�[��rl���ڮ�
$�q��P�ϵ����ñ*���f��>
��|�%��ܒV^��P$�6�pv�A��'�!J��oz�6 K�!7Vj1��ƛ�t*:�[�T-Ǡ��׍�B��w����zO-��OJ�}�,��z�L�Tq覆�aC�g�ݒ���X���l�鯁r��7��1q��" C��Z�I&q=@�+MO�H�u���M���CoG���A�� ��g\n,����_�����(���w��]T�k6��dc�qƶ��<B$S5q�pّ>EГo���4gja�aDݖ���>to�_<��$5JgM�N����G���b6�pѣIO��5�)��%l⟳�?�/��*�k�!�����Rkſ�W��h/[��6,��-��3���0|fNԮ��� ���k}��K�c��J�'rW�R�T��K�N`��/#����V�!Vw�-տ�u�=�5�����L��5�%m92��)%�+�u������- f��S"����%�t-a$ȒLŝ(�`jec��$^P��������|�!r�_��?��da���ۯ��j_Q{fy��"�~H���4�]�������J�{Ժ����w{�CQ]�2i*��f��(��򣽠��S�(X��)V��h���k���
@�[���%O��ɮ�U�-�13&��,?��ĒO�����e�%ݬ/�����˙a��7,1#c\��Ϫ�\���%��4�p�o"�ģ�k���ؾ4���:5�.�R9�5�f�6�s���z���OS�SX�Ԍ��(�0D'H�I8��{\U��EІx��x8��|�Q�U��7�b�"�h$M���)��wQ��L��'�- 2g&��o<���"�-�=A��������)�7ʲ%��$��~�C��7��/5mG�T�W���芆Ȁz(�Kʻ��Ȏ���:&E�PR�IgS\!7������D�@�>��\	�12{��gK�������yz�B��¶�'W�H,����=-L���-3a�b^v�81�����;Lbx�;^	O~��q>��j4�|�|��g�wM|½r??.�tv��z�ߏ���RV� ��S�M�_|��:�dLX4�B�u5ّ`�����u�-�ChB��j�*�4>jj��.0�۬�0���f�Cr����1��w�j��?��<���"�����r$�# ��v���-%YZ�KZ]�$�"��o{�C�'��})��Ys/j
���}x�����YǢ���7WD�s��X��R}���y��V �y�^۞t&����� _s��$��]�}��I�"��X6A�.�2/���--�&�Pb
��|1+;���_LW�*LT��D�Ǯ����Y��f����W�ϝ=�Ƨ�E��k�K���T���������{a{�پC�>����	��U\��R,'��ٕ�[�`0Jʄ�1�>��h"�lP��a�n��F�K}�x��#�%paT��Cx����K=��Ѝ��JK����xFÜ�w��7�A�=7�FE�op�Z�m��T�NW
Bk`�ڎ��*����-��@Mؿ�7�bw���+�d�O�|U�rj��t�pn��C �>4y������835mS��r��_���#����(�#�9ؗ#���^syR���|����B�y;��63ς�;��S��L2�^�v"6!��A"�����b�d�h�;�d|��g��>-����+�\D�a"����ӊ�[�����8�@��ǔtK��-HI�w�kHK9��? U���9�B@]�U9c��m8i�!�=��H�����şz�f-���X�upVu��9Ozj�N���
;~����:4�*�=�}�u�~
�=.��d�@"_U���&7���>Vl�S�p���PM��.�*�V~W麃�5�C�@����ws�iA�-�jY�����xf�\b�����U��Qי#=c�P:�uxW��_^ [ƌ���E|�r7ufR�:[��ln>		�!�I�eYL�����{2�5z|2���d77���	���ō<=�2��a�:~:����F���V�݊*Jb7���_�0������Y}��p���z����m箚Ʉ�����B�ia�CPE����袏�h{D��h��!7I�~�8&�i�v+��1�D �� n?n��!E�O��uڅ�,�P�&�,c�k(�]z�l�,�}3����9��"4,���b���z]u��Fjxsa�Q
��� ��~<c%��ꙺ����E����D<��<�k��8T�J�9f�����5�{���z~U��$G��RQS�^���K����^��3nod�r�\?�V8,����`y�V����Z��a=��$ (�thr.�KE�-=U1�?��ׯ��Kڸ#4�<���~���ȨW4�ßh��Ĕnj��L���9z�dU��.�C�rg��`Iy$����-���~����z�r������(V�4�ߝ�é7#��iV]4$o���"�f]4�s@��3��Cۉ�J4U>�g��7ț��Q�"�2r�p�&*��]BSS��ا�l⢨���|)���g�>ܻ�ԉX��H���賃�����w����	�$\�*>���3���$c���N_��������c�#$�E� �� ��ˤb�MYD���6���.�^B�A��|+��Ϋ��}��8�[uv� 51��!�����p� ���"e�5�p�O9KC ��.�h��@��L��VÍ��P)h�aq��9Nj	CQV�5B����P$�I3c�^��fc�v'V�I�<~Y&F�$��F~K3ubs��b�;�r�H��1�n�XTb5��`j�kz��ګ1��6�_w�m�E�j-x���v�b+nU�ȏ�ȕ�,�\��$�.R����xj�Z_ �g����Bς8-�HOH�w�LǝȝY�0�����9ui��S������jV���@F�%��k��a��)] �Lݔ�C�O<�Nǎ�\��&��3I��!�ʔm]"�,�
9 >��nB�Z,8��rV��' !Nx���&��(��`h'���)z̀�d@�ӏ���R2D�4���+��	���DO������ײ�>i��"M|4�-���'7v�%�n<
��Ǌ��\�L�*.�mk�>H����*Ϫc�*R}����1���A̖6���N����w�+�3x�R���$(NN�kdB�}�A�l�I�b�H�]9w�e�K�o~IMs��7�3�:7�������p���r������d���-۝�����-�1�@�7�1�Kz�����4	5;vh�5�7��O�7\�p�5���Z�]�E!������)v�i1�ێ��Q�C̦ ���L��*2'4�Zdۨ41?6�A���yIcbC_���8�6�52����LX0����|���+b@H�e\�@��ާ���]O����&򺀃��G;YE嬆�::X��bڤc�c����������Գ' ��.�.y�)�����b�>6p�6E��u<�gEKCD�۫:!su������,O�a���tkB�`JY`��Q�{���D:�"q�l�'����$E�V�mf�H���	j/$`�_E�[%���8����#��������&��d����΢�;?1X���5�����Le�5�pe8_b��}�w��ħ��Ȃ֝�H����s���G�B�r��:������CKY��սWw�ǉ�.t a�����^��O<V]���.]�1�G<�r���������-���I2}ʴE��M���z]��3ԛ� �Xzӭ�y!�K!�\�2�t�~ດ��7�4�GM���T��;����n�g�~��:�4r8�F��CcȨj/ XF�oG�VCP�)�;���9C��ߍ �բ����!5�\������"��h��Ѷ�ͪKS�)eS��� >9d�<���+��y��,�mLA�)�x��&�1�7D%�wl�K�����c⋉�F�=��0@����1����}���j�äƪ�ًn�"���٥�60�%s�������渹����o'��HT�=ö_ӕ+�4Ҟw�w��n�/��z���%E��/A�E??�]|j����z�,-s-'&���+(l�����r,�$ğ$O�6p@'[y��-('ȨY��T�N;�Ԩ|&x`1�$�:O��hLnYbƤ��`����S9&l��P�)ė5�mi�[�u4�	AbJ�_���v�:$߁���( ��������j�_Y5|惂S�x��{��c|SgZ�P�a�1���.�6sgqB��1�x����	��i�I�{J&�=�l�ځ�H�Mn� {��2Ktеw�d���a�tt�V��Pyaj�#�>�!Ҽ���]�`q��}�������饉w˹�7U'>s�'{�}
8a�����*Q,s<�۷�I��Y�:68�9���
UB�ިac�=p��Ȍs���� ��|F4%�m���i?��S����A3Ϗ02'sX�=�-J���44��(
2��kX��dbc٬�#h�XQQ�D��,Y���(T|۫�ޑ��w��§�c��$[�jnZ��<��Mj�ϯ��	�m��=���Q��WЦ_ws7�V)`Ld0��w�4ȸ���:��u$<!#Էjj�t�sş�������\���NQ��t�o��K���HL��E��`C��A��������b���o_��t麇hsv^������<3�`�ܳ�f���^�8 v~��{厗v�S�Za37�H�����]�7��2�w@{P��8Z1��}` � �!2s�çD�<_j�yE��\��(S�2���
	5�9_ͱUj�!�{���v�z�^�,:� ��	ssEn�D�[��S�-��D=������Qf2|��&�(5`�e�Z��"1����0p�97�S� ��c�R�����AC�yl?�K����E��PK����ٛ���O�~�2����FIX�k���h��7/I;�I��n��@�������D"H��T�2j�	jOY�K�����m��{�rc[���c'�IZJ1��/�s�{	�� ��i5<�h�YZ�?W�4�eɎ�C�S5݅��j�
8Ue�������w�r�H�~�����ة�8^x���V�/f�n����9��fm�/=��]��U]��W���1Ig��6Пˮ2�E{����Z��S#hRv ��E�}2�@]M�f&.�s�M~��ޞٗ������-	kO2�-7�Ƚ����^R�Q�;Y���рz�E��8�G%��V�؝�,y�Po���[�9���&(~ēd��ģ�so\���L��\ ��ޚ�v����Ω�V�h;��Fb1p�t�-�'��a�8F�@U_��+����L���i`þ]���ٚ80B��m4��m*�ݖ�NW#�4�w;L�,ף���0ݯ�C��q-�&i#�8��@�TO��\�#��.KU�E�Y�L��jM��$X�jS��y�]�� �"PR�#/\�Q�~�Ye���|���C/C�480u��q$�v+�Q�ee��/��n�݌=|`I���GB��)#�T�f��סD	�! Dz:DEbnŜ�E��q#�v�C�=4~� 
1ʝق����V)6�e�7}*&�&���t�\c�Omy"}JM���H�&�R���Q�)��
dl��1����,�N<��$ɓϺ�*n臢o��q�
�P�[p���A�:'	����kd 6�:묄�� T�����Dw����i���oE�}49bP�i���r�O��`l��b�,� E�kd��T�6ļ�]
x�Rc׌�s��lq&;}c�����{&?�<�r�@��ȎL0����/xz�� v��ѬS ����s�L1�;�
x8Ď��۾�wJ�#�l_՟�\�*ۿ��r��,�Zm�����|ǷY�>����(Z�va�J��������+LOT^��&�k� �o8K�(��R>|j��X�ܪ}�I��Q�i�1:S�/���Kc�sSnM�-�8�]�{��_Uե�g��pn��Έ�`j���)_����Ͱ��6!�U���H^�V��I2�+���vdk�?�'f����>o[p;�B�F#s�"�G�1NMb-�]_+O�̾���X���E� ��P[k��9UY-�HU����+��@	S�v�j)GQ�Q��*B�`Wd�"�@٫�K`��no���+��dď9�r	Vg!EY|E�L�o[ʷJq.�"��S2��.>d
L���7�ݝ ���R�
nn��t�Q��w��'���r·~ҶL��	UD��D{M�����S�X�����3[U0���!��^���oی9�g���1�Kph��5��A�k��p���i�d����ty�i���n���=�12��w���� �4�q�	`��SI�<��j�j��k0�O�#9�Y��`_v\)�n��y�;���5�|�X��:'hL�U&�t;{�]�y���m�m���Ly6�uA���CeS��Q������i��z�(K{S�>:e�
�H���ۄ��qf��ڻ�]'�F�����?t�ߑY&3��f78H����x�gX�,܌�ؾ����j�U�~M|����'$: �D�جk.f�]عx�i�Qre%߈�j�����k=�Be�GV�LG��`�9����^:&�@�UZO��@s%�����1���!�*Ɵ�/���@?Tۈ�%\��oq&z����C��+ɑ�� p#7��d�K�k� bM!?c�m��iX���;%����#!w��R�!΢�a���X�C��䜇�l�p+f 4�+�������\����;�w���<:2%���S¤�k�������v�
x2eV��9	�>`F���ޕEiջ��H)����I�9�������5
ۼ3c��h�j�EfZ��؅}���A�W �P�n w�,4_ox�M�ww�Vl�[����fd\{��F�>��P9xk�Ka�p���
A�A����,�=NL�~������T�J�� ��<E6f��6�r�����>�@w�F�f���R�w�Q[<�م�\W�;��WbV�r�F��AN���'f���t�0:���u-U�b���!}^����D��ZM�aC���;� 5s�"����wnـtw��I>��6Ѐ�k�onTm����(À��[4��굲�(Ѥ/^gdZ��9�m�.a���xN9�ޤ(���U�CV;��5���&^��4w'�NQ�z����hl�E\cf�s*�n�L��On.gdM�!���{��$��|G�R�Y�*��'��DCl�kCr������|��4Pa��Y�f����
ip�!J_��B�`�'=lo0R���~Rѡ�n�	�~�,���Y�J.kcT���P�~ �z��g3-�4���<���&��3�tfܞw��S �x�\ᵖ�%���#��z*��.��:?���qہu�JW��	�F��M5���s�		�2 8�~p�����>�����關�6�茱�C�%�~.�/�	���ڨrP�J�1R5�_:�����9�
����f�@g�?��6���OW,7 ���w����}-Lq�¥��qQ�����SMhfE�����}�u��j=���f>��0E�0+��Ͳ��*S��í�?sW�3f���1���b�p�1�0)[EZ�m�cǰ��RiBb�u7:�����u��x�;�a��&���PR�$�/(��"�F
�ʼ�F�	�RS+u�j�9��G�A�<z��&M(� ,:]�俽�Ƅl�w���ζiwj�\�fu�
�	��*r����5m��B�S�*`���{2���(�H؏&ާ�@I��ȴDK5��[H&�Q�R�.����ы�Pf ���H^7�c��#��74ɞR��si�p�O7�+����Ma�pBpҢ7hB�	���ec$��L���fu_��U5`��}��y����)TMO�^��|�"���/t	�P7~d��=�B�<����q���[�xw0PZ� �|�m�H�Y���󫅗�fZiFU�f�vQ�Q	-;����(��N���/�,��@T��|D���I�n�hW���L���gD{��&���~�8�b]w��L�}��|TÙ��ML�XY�G;��70�E��½3�X�F|�F����#\_�楶��|U�7���^"(P>Y��?XU/�^������/��u�̧Wz�;�) �g%�.��҆w�2�K2�~�,�k�I��2Бf��fB<�;=��	����_�л*�ߐ$-;��l��պGE|Frs� �a���EG���$�+��ºC��rBl~��K��HuC$H)���h�-?�L���c����l
i�rb[	����0��T���2�_4omwJ;̄ �lW��2���	��y�������4뎭޲.j�-s<{D9��*As�</ݭЫ#�0N�J�irH@҈�W&�,��g���*5���pP�>hՃƟ�^3��G�����φ�>��b�I�{Z��Du!*a��f���J��[nE�ODŷ}�wS_
Po��h�$wq��d�c�Hm����b��	��J�48�͛��1�(��"8P�xD)s.���'u�D�q��-n�� ��ͺ|E閘�&N?{ߌ���/�KGd���/��/��xP�`!����V�e��@9~bg�Z3P��PjL��=¶��	�,u>���ײ:� ��B:�G�,�zg�:������܊Y�R2}�>�]���ЬxB�zl�Y+3ۙ�g���RGJ
�8�)�׹���B�e�]�s�D��1��Z>�˘�F鹧M4�\�������ty�'ܤ"b��<Q�;4*��5�YXI��D[Pu2�\PYү�i)��w��@��v��;}�=�բ̸������b���KۅrL����8�ʆ*O�rc���) ��&�yx�&[��s���޹� �����'h	Y��w50/u��!\KF�G�i	��=s���x�:)i�Z�k�Oҋ �Ӧ�� �O��"W�\��=u}ߔ�r���x�ݕ�e,�ηޥ\����u�lo�����[B���{!m,$ڍ�}���(䕾���Lq�b��&��д��1R��5p�{9����A"E͗���E?=;XZ�{��7*O��6B�;�l���3!^�r��9��Nyo=B��n!����� �#��_>��/D���)�㌊�j!�u��d�BH�QRweY�����ҳ���}�K}{�#A��{��M6�6�ۿ��RE�po��C���tf��B��Ȕ*vSv�s*�(�L�a +=V�W��*��]=�ib��������Ҩ��a���Ѣ�In��5��&J�ߥ�1,ы:����=� =-�BA�����z7
�m��.��k
u�m��g���ˡ�'L30���������?MV4�:�,���W����
��F��z8�@+�p� �Zt�G�ޫ���;&ڼ��g[3�3_	ʈ����t/�jWͩ�6��'����n�6��E
���B�Z�k�t�؍mUA��~��sC*���<4�\�L,꒲�R�JO_���wz���@��F#	J�F�����J��Z̈́'��Xc�]��I��KQ�z��cUP��r����8�+d�,�~����n�KH옴b�y���f�\�a��d�(0����J˒G�H#p�¢����`�" ��F]x��ys�����PD����<|?��܌;�-�%8^�29YA���J3�O�:G,�w�hzf�ɺ����v�=��`c.�EM���Ub�x�p5�.��@�c�֥��ǋ^��v� h������n|�a�E|�G����J��R��*0��w(�����;L�*k�ġ9_d�߰c�#娖�x]8��Hj��r��	7j[����Irϡ���M�!�)# U�h2��j?AL���?�i��W��W��&�4c���_��³��H�7�TA��gS\闘�����m�g���c8�-��{Q��jCy�3��\WNJ����G�����v�s�7)�� �0��4��h��3b��6��Yy%�b<���19�.��q?�<��P @��Ւ�
�0� a}�����yiPP6h/b�حD���Lc�z���	r1zM?�V���|�*�M�>�*�d��}4�Uj6fj%�`	���� ��ݣ����Z5�����Z_
6qK}!���G�Z�8`v�n2����̧!,��V�99UW��3��{e�8)L��� �H���(>Pmw��9ో髼�$D�(�G_wY����?h3F�Vi�A��'�,a����C�tN�%H�Gm
�"��p�g�+	ȝ��7Eؐ��΀8��7I��2��&U�����3|{a�=����{���|\���lW�9Uq\ѦSq�t�ñ�9%+��{{O��J�T&�oXb��ʃ�Б%��NKO�_��a�D ��	���K�ޱbu��K�>����+�k��XUl������͛v��<W*|����f)�8Б�<ȴ~���
�ӷfK?���Ѱ��ur�\�2�����9���/�NQ��z���p ����x�|�$��Ā��8\,	�ڍz <��(1���7���H�X���>��8���ؗ��}A��/�P$n�[w��J�RM�$m0J;�5Y /vuϭ��i����E,"��r�����6y�0N;�����¡*;sԹT�4s��;�"�z�Q�I�*f<|eY�s�G��p'��4�A&��Py�-�q�E����<��k���\�t�l�6���cp��|�d4��A���K� ?����R��꠨`�c�K�*}6���v�-�F��l�t��18�}���>�r �0�;s�����K���%.�ԯ� ��ki'�ѷ��1�>���C�8�Õ�#Q-�gS܆��t�g�̈)HQ�����b䎿�)�t�-�ŀ;�n@��6��?�Z�%ars�(Dz�3E>O�!Hɥ"StFs�$:@⡌#D.
�;<_�s�|KJs�b�?$y@ �0��-����H^a�8,ơ��:�㟙8�	���	+�&����i��#�m19i�x�[]��L)�"+�X�☍b�:����+���o=�����b��Wp\�߉�ՏP+7��yF3���2���L��W(�Z���Cǐ���>�PB��Pטf0���D�L�xR'�0I7��z��<Me��?��̂�n�"'�q�@	�8e3�&�m/ʞ7�<�+� ��k��K]���䭧#�Bc��&	.:��@� �톷��,�Җ⍷a�������-��i���|}�*������.�����]~yې\7}
F�G����"����v�4��P�e�=	�vE�~�)�\w��˰��o����]:��g �:M1�����<��Q�aG�|є�:�H���$�9�{���N���XFP���h�a�͚���T��U��� �]Ѭ�kQ6��oˤ�Vb��F��%�+I�Z�"���2^���&�Sp���HU��h��l`�T����.�`�-�P����P�z��d8�ᵖ�`��x�ݱ
��H?����0+2Sk�]����s�NXS٬�B�-[&�R�	��8�@: dt�$�o�������)a�e�9�\U�������TjM���6�5ㆄ{n�B;�z8�օK�,�������$"р���83���)U}���T�o\LB���h疼[[�e�1,Z��vL={t��Y+���\"��]'l�?U�bR����}����S�]�3��y@.S?;n;ߡJ��ZCJ���m���/'GQ^;?���Sݗ�8һv4.�'щ��x_���dԟV!��6�s�}��}��x�}���7̤Ŝ�vs�i��Z�^MyIP�4+<g'�FH�P���i�"vd*���*����`���)�LI��9w��f�6�;�d'v�km��I'�_��B �>�Ǻl�)�48k:��(:� �GmBC#X� (�S���z�@{�Q�'����8�̌T#,d��otޠ��w�⪍�_��G5�p�;L��9L@�Js��%�像&{0G�X��,�-h	%%s��p��f�!a�p�2�k4wB�r<��A����<���h��F�\ҏXq$I�u���;�Z�d�<^_j�Z�ۏ�Ĳy�m�w)�,�E�.�������k.8�8;������Ȁw�$*��8�ʏ���>��Z����=?M~��Y��]\d�H�����i�H�2;Wz���T�Qx���~uS�TOq!V���-��R��P��o��:R`�7{ć�4�mp��ּS����k��1�����9�}�}T��I �ȹ����(B�������P�]#w �]�w�]v�	���H��԰��
����T2a�W#U��>��fD�q���<(�x;K@(bo��jR^�gM5�~J�^�qV=��ȍ��ёf�0}Edo�n�x�M��(�O��::rMH���fޒ6-�!�鼧����.V��М	��jˢ���3qL.P��=|՛��p3,�;n�40#لZSAM`�꜎y�a�����ѶȌ�l��a��|�0��4�)iq�^���t� ���O���t��u�D���=�m