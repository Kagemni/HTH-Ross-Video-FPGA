��/  �F�o�~���W׊�m0�i�14w��9�@|�L2x�����%ן=�M�,�d���g�$���-�y{#mf�D��T\M�Cޙ>�X�룽�Q�TRJG,O�w�/ۣ
��x�Ӵe�q� ���5v�����hz���>6� +�9Yᢖ{k'BE!�(��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�UtOU�0:{j�IT���]�g2�[
Vf3�����=���у6)�R�@���k�mBP��xu���f_���1]%�sp;Cz�����D��t ��D�DX���ל�+xk�mH���U����Utʾ���(��+��o&�tUf=�+@�D��Y1��W�<2��f+q~��Ƈ��R\/u�2���ʓ���E�Fs���{<�`7ݹ$=y#ܧg�$���i>f�*>Zk&��7�\�ܰ���_��G]�y�U�7�S����yM�Kfbf���l�ܮ~EYj���y���ʤm��܅V���B�N7
�πM���{��k5��.��.Lc4m����80�@C�{��zۺW<x�QK��?�;I��3vΜ�*�~����s{72������>�~��yW�JM��cfҪ[	���O��Z��A��m���	��I�.�ҹ�7��S[���}���)0�Q�E۱X�	��_e ��aB�<J�B�/F����
�:�ri`�|���3z�B�l�f���a���f1��dٝgV�sx��W�/ʞ��IY��J�!=B����S���T�8^�w֙�x�� 7�8P�A���x	��e2a�Y\ӎ�wy|B/�:���~��	���Yغ�[xg;�
p�+�g�ʢ��OG><�xx���,��_�Ļ���SSN4��8^�2���7+��50Xjep�*,w�u�1B��%,��������p]��}c2�������,��,��y�<��;�-tq�Z67A��5Hp1>�a\v^�� )E��ra�x,��l;&Ԭ���1�����΍#��c��bޕ��C�\�˙{-�`9��LU�qfZ �瑃�� �g�cr�����{k��t%�tI<����1Z�!ߌ���.5`�i��2.9�>k�I��{��`�JO_T� mq�^����z �����N*�nf�_�d��T�[�W�?s���ҟ�X���2)n�ާ�am��-�X^�@��ޘ���=�~ ����i*x��S�Ǚx���N�E�#��PLu�{jv��Q�&D���·Q��p���X3`�⣹����&��:&���3v���L�}�x�c�`q�%��BY�D�*�f�S�L3�b�A�Y˕�4�a�B�'V�r)�e��m��n������5�O`=Z��F� ����n�]��R(���Qm�P��20��o,�`�q�x���7��WާX]Iƪ����t�fӣ��5{���y��`Գ(�Xb��;)>���=���J�6n(���fXԕ�1D^n�� �w����)rs�t-p"�@I ����l�fj��#;�c�<�vMn<�O>,�zlxWI�B:/Eer�A�!�o2�n��@+⡟;5M���x���r�h�d�}{��)(qHeX�����H����(1=��I��ŋ&�#g#��Q}��p�����~���{���Z+Sb�9d�O�Ԍ�ŬU@I�z��(��C=v��>dk�9�|��5�;ʜ���{��~V���\��@�yp�0cJU�K�S��-��kJ�!�*��.H�HG�oؔ�{>6�L���f�(�$0.�.�J�!�E��C�(��VvU�Q�J�a�F]`�<@M=t�e�BqqO�Y}Z��i�u��V�{�w�x��L��yT(�\.k�೮nu��&�m f�V�n<��+�����j�IU�9�%�U{��h���+���H�K��qw	��.�Ψ�DӤ� 8|	$o��yD���y蕩A�;S�&��.*����hq�Ṇ�,}|��/��j�g�r��p��r�P%F�� N�e�AA&$A�E�e��>'�M�+����\N����b��:�2�lZa�k�3�f�M�*����٭1�[{�OG�G5xo'�Y���N!�9�\��Z�G�&��}��_�T��B�G�������߮�����?���A��)p��� �����IY����)Nxʣ�le#��;@/�_p�\O�±�����8���!�Lx��� 2�Hi�"�K���:s�l�x��Y�?toq�K��FZʩu��fV���RϤ��3�(鼚��ځ�oD�>�i���Wf����(s�{~W���e�j�#��>F���RJ��YJ(��4���"	����ۓ�5E�R�hN��W��7(�V�b)�U����3�B�aV�E�7�"�_��.31�m��`��3���_͍	Y���X�6��ˢ�a����T����9�L�jZd�L[���[�׫,���E��u[1�#Z�I��u՘��dK�d�G�&j���d*�������z��l�С@�X�GJf<˔�Zp������x݀�f>��	[�-Oc�D{eR^�(w?��T)1��d��>������&]�����`;6����RY�ya$JQ,�OH��JK��sX5ʰl���s��_�v�M�h Iu����͚[J�X�$��0�^˹y�2�N}ˌ�3��h�W����Iw-๜�I�/f�i��ox>�BiK�ai"H�1�V�[�4~��5� �7V���JK\��49T�M��W4ҋ_�S��c��-�+x���	��[�D˔&�lR�������5p�>}��x�Ij�R�4<�2KCy1P�ֶ<yfߴ}�8Ă�HLCQe�r%�
'��u�#C�����>�]Q��g���\�҂�h�)}����P����rbnA��I�B�NZ�I`Jq�(�W8R�akշ^�;�G�֓RW�͍��� �@�x%%�si�LO�J�>� }b��иْa���h-��R��V���mre�<���Ľ��EJ���O�n����6��U�`A�\��&I�u������Q�	�g��e��#�yD������쉑��8������u���i���jZe�ЋqN�~�iQ��J�/>Qٖ��J$ �ii!` Zĕ�� �=<��F�f=��%m�9��D9��~f�-n�P���x������-:��E_f{]����=������efe���L�O݊g�4��}�%�c�h �Q(�����ժ#77�c��sPPA�������'t���A�b��)�D�����g�>Ȭ_�%rwEo�S?�D%�o4�iܜ�G"�0]���p��ݦ�D��s}h�.R;�x+��� iME%Z�A��U�®�e[��R;�y����ޗGbuwgp����?�;<��"�]$mz,���$W��g��Sl�"j�<�FWٚ}g%�Y꺗2L��'"��O���Yk�wqu�iLc9]�! ��͵�¹�F==q��=ߧ��{K˝�H]�<1_��6���$��GB��2��,w��gUj5��m�~~��֥�����;R^����[�|F�R�69\�%�|��yG���y�H��ݛ�9H�����b�M��N+p��s�����O�z䰄�P�	��J9�a��@TѮ��E�!�[��	vY���͕��IEkU=��vy�YzG�эd?��H��g��L4>1�:O��\PDj�tƹ%��p��~?��qv0���K�,�	����>E��������MX)��Mtt�(7+q!���eD���?�� �)\Ԃ�pP�P0�>���7X`�J>Yc@��7��њS���K8@']�q��͢/.(�
�1�U_�X�8Ml���EC��l�п'���G��c�p�J��C)��X�ճ��1&��e�݌4�i"z�:󪇨��2-�b��vP@����'UZ�L@��R��A����e�h�w!��ٶ�B���8�c�$�E⦤�W7x�ʜtG� ����!��قM޼WM룯���C��"I�}�}2�Hi�tG��.c��w���]���}XS��5M�v���}pfAwG����j|_�5��H�k.®���%�?����Z�K���)}��p�Ka�jVM/V.���1�
��`v�I���;Γ�ݽ��x�,�H�R��9���Ag���ھ6��پa�[�c�LP�c����M~D��Ǜ�Q:p�0ŁQ���h�!��VP��W���ͷ��},\�����"����b�چ�H��?}�M��Y/w���|�7Mo�L������FĔUuH��q�������H�ֆ���c��ӑMZ�Y��h�`� 2�vC�;Kո6�SK�[����&��j,ӠL�ǼV�Il�ǰ����M3ٴǷ��e��8)1�J���ϗ���"(i��Y�����YR����;07�)��$%����z��'��~?CY&�b�6g"��4�%��;{��u�AO~D�1xDwE8��Z���<�-�;?pYX�e-AS/��%707$��a��K���}#E���;
���P	�-��͌c�%������v�#��Q�X�<�紧�$�_0�|���M��c�p����X�J�ȏl2��'�N���<
����%*W��U�ȆE��M_8m�m�g���ԭ_��a�Y�K��g�|�N�zY`�-T��)Gh-є�?��3��W�����<����0R�}�`:�Jc���2��u���Z�>I�7���Y��A���#MS`j��ol8��k��5aȟJc�bƕ|q���HώE؋L���q��^��:^t0TCS�ӫ��F&_g12`͎a�p���~�Í�@k��Tz/2�D�/&kQ���w./ʳs��7h�Ъ8G���t��@Tv�$cW���P]t�Ej0�Iv��)���sf�D<M��(*-�]�g�7��𧓃���X�� @h�Vxݴ�F���*a$"��.��ƨ�mD�e�uޔ����?J�����
R�4[[;�0y4ߊ�A�a�(YbMݸ���0����F��k�T�$j���mU��,� c�c:���N9h�DFt�����1�AL�҈�@��$�x�5�}�YxC4�bӓ�@׋3b�ǇW{7���1��馀ޫmf����S%&��e��(�Yq	���l��]��ZC��}��ܧ#��˔4[ŪC���y�5J���OXv�8K�� �e�qĴ��`����M;Hf?�xGC ���#��Y�p|{���I@�W?�fM
�q�`S�2;��
M�mk����F��k0�)8F�R�	�sp:~�N�KrLj�"�b�^7f�3*�Ir��=V�R�>���
rR3�`Ó@>=�Z�Xw����$��=K%��:Q4&�+�60/0h�&����: �t��&S�.�^s�)��C|-��6�Щ��v{�i��X"�}*��c�5�fn���� ˚Ӡf�!z]/[�B�y���.u��PJ���8���h|�M]��S�u̢�'�����c�,���*_��S��7�#���>��E���)0'��X֦�%)%z�e �[[n�s�����Be�В�j6�{U��pRic���f�D='����A�;��a��WcG>�c��E,�L�A���xІ)���'r�' ߤ�ee��t 2,u$mX��m&���2��h5�c���^;Wκ	�}��G��`+�[����Y�G�9���:X��y�d�0�Њp��w�P������dqa!�d������7r�u���C'f�	����b0ꦷ�s�g�
�$:�h'�7Q�k���O�Ӎ{{�x_޸_V]����Fk+��� 5��$,ɧ�����ڇUJȳ�Hs�����Թ
��_�I.����qNi�R�篐�ɵ8\���g	�I�z��l�*��Og$�e��z����Ӳ����`� ��m	@�CІ�lG���غ�79�<�	��R��".A%��v�7���Vnc�vN��PbR'��np��������
a]Y(,��5�۠&�҄%�P�Z|��l��=�?�P7L�D��M[ef7����K��Rf�7.�<��w#���δJ��_��bu#�o�с��|���l��b)9��S�K+���+���%�� 7�o�FhT�0���"�r���q�~� ��I�ڽ�i�c4����V�x%�����~e��֓2�L��0�{����(�w�p�?���}/���KB-R�������cңlf0��$q߭�;m!KVEtq�^�{��6�q�e܏z�N#�gd#�15=�+ ��	c'e&���b6��1& �U��Y��.��fQ�xG�m��
�[Q��y� ������NL.m�`>y��u]�8+���Q>|�1|�#�ֆ�C !7�WV���RH�8O�J�F��9$�M@o'�����7DA�D���,�Άq��W��ʍe1��%��&�'�u�3oMD,�m������?��̒)���z۸[�w?�զ���(�q�����<���l*���t7=gA�u�<豌�D�:[h's�v��t��h��U�}0��]�)(n�]��2���Gt�'m��/���}*v��Y"��;ě+N�[�v(�h]�w��n�F^��9dn��=�Uqtl���_�yb��3��I�_s��(�QZ/����FOxT�f�7�G��dg���ԟ&j��PD�������w��(j��ܷ1E�~��x̌��q��PĔٷn�k��6�Dj��C�v�B�s!�OS= 0'(�~����%�q9Qt��I���~����w�����U/����2;�c�`Y�r~��Y�Ĭ�C���><q��V?!g����V�P��%�;�-Nzv�n�gذFB«�߼
D���?xb�#��SK� H�*��)�$*�8�l�(?6IF��X����#����x
s��L�{�Z)a �PK|��Ķ/�%uP*z���k�wbQ�WV�u�6���&-�3j��A�+
0,��C�sEN�r�9������t)"�J�\���F����c���:r�����E{��H���;��>F��9�@T4�5�����Yr�p�r٠��MM�Z�3��I�
��o�i���a~����NE����D6�Vc��	}P#υ�����	x�.ޟ�J��[�c���P�8�C��2�?�sa� P+�(�F��cN Gk5p˴�2�sh1��j����aZd,�u���WKC
�o�dT�M��Xm�󎸷f��Gb��K ��Da@'��{W����މ�h��!uk��|$��8�{���tB�6�z����c5h�������P�H��Ú�� �F�CY�D���̮ߝ��<�<��ue6א�p�A�(�s4�����_����"�^=u���$%�ǐ��xnŉq�O�aJ-ʜ�~DfI(���d������٩��|��_ω]LU ��Oz3�`?���r�rL r2�T�;���G�q��4p���G"`��c��������gA6Ҿ��I�`aV5Z�]���j>�����.3] NH�vf��tș�����l�:��PU��n�\Ӫ ����Ļ#qb�F�f�T�8-#�=��"���ʭבN�LXB:Q˖���C�_ {�.	ɿ��d���Z�F��c_qaCzޫ)v0`�!�����\�OT��i%���[n�bc��_�c�_Ny�r#y��'���խn.�eݍ��Z���ۨZ��cM���G&N�'��_����e���Bz�-�B	K�$$��4�A���htVe����B{\�����5H�~��Z�^?eP�<o��J��W+�Γo