��/  �9�X�[k�5��j:W\���(�Qq���\�6Z��iw���2n�oҴ��)B��.ƒ�S0����\%���j}��#La��I	;~�k�[~)����AG�"8B�}������L 4J���R5�e�w� w�	�&�vs"��LD�3ǈ�j.��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n����~�@ԁ�du���C�""?1d�2�?:������G� Y@�p�m��Wى阠>���AIR�r�n��"Z���&?�ۻ;����C0����%'�Yu����S�֑7��W��~<�II�����U��2���5�>��l���D�~mד+�����?4c&h���T���y�2��\9Ǫ"���o*��o���y�*,�)�/��bFDe(�Z ͨ�5�O����h�؃��(;!ь��Y�e�13 ���ޱ�Ǐ�7ʉ�6\,V���@���l���7=�iN0CR`�&p,-���8�Ik�3Fl��ղ����4�>����?R6��0�����j���y��WD��5�k�J; z��;���3��hټ���� �O,��w��:��j�a�[��Q��2����jҍ�VQWѸ�m��ѷ��i٣[Nc��c����9n�+��E���3A�|4��N央�"�A�,��y�%��J��Y*�ժ~O�EAOFL��An��"��E�����(����$��ps��k45�]R�N�Q�ģw�]f���=��楘��L��h��E�19ɧX)�<!fUv���ճ%%��.L�z�Z���{iqJ���D��5����!٩eq�8B���s��6^5)UN)��F��3Wc�,�ͿMw#I{���6ד,G��F��7�%Л��)�C8c�`�<'h.�}��7�\H�򂿧
>fTW��0j؊GبO^�^������^��V���J��&b���)�b@n�`}����e9��m���/'g��[<6�SK�D��6��u|����=���L9J.�`_�)@�����gRk[���cb{>
��;�qA���<��Ľ�-��n��ک/`�0;~l�@��~�X����	1��v̽���Ă-p���Q;V�t�վ��A�Q�ņx�®��}Yx�*�i���uL�f�P�k�.?A��ǫS.BX����Ӭ�[�]��fs�)����酴�� 4֌����f� z��o�wz^����4��T:8��ߢ�Go��&f�Á�v�ߵu4۾�|4��c�sN�M��Mj���r	��ݎ�TD���4�%/dc#��S���]�'�:�n�C�.sY�RG��ȗw�[��kh��^{s��YoQ��M#�s�{�B��/�<*��a8���і;�탬��~B�j�`�=��+���l�}�Ĝ�`y�	�"�)8��_�~�Gc'
�4��l[X����Z��$g�=L> �G�������h��9Ѻ�Ձ�r\���'�B�Z��2�"=g�2��3&�eO �bN�ț�4���p$�X��&q�/��p�X�c��Ç6�S�P��3�����R�SP]XJP�\ C�QM�B��@Zd�ѺW��/M*�/o	Y�I���4SK^��df �a��a�:FO$C] rq��3	N�h)���F�%��ƗJ�V�+�M�^٭�+aZ>�HGX1�x�Y﹎��Jg�R������ �������������J��`��{
X�Il�X�Jq:í�Kd�*��f*W F۪�s�V������ j�^�W�n��:U�.��?aڮc��i
a�U�����?�]l�∌�GS8c��Xq�u��9<�W�^��= �߅4E�d_p�|�œ�*'�d>չ��>�U�6-Ϣ�8{_��gE��@����,.�M��^����eyRx�FX?����0���&�#�7 j�/<1D�%Xe��Jgc���R֭���)�h=��s�󰜮Yj;�V.��F�L�]�Md�kEwU-]$0�H�!�Vd+�%��Z@��Sr���,�q?x.��9��_ig��9�]���Y)/��!�\"Ҳ�Hn�*邈�� ����	���-;G����[������zy����<�3��3
��WC[��- ������/P�A�[���8����):Ro�7k�q:�G��y*~�E;{�aa�$�DY���A��u<-�0a,ǇC�y�n�����>�f����
���6�.�I���JA�_q���g�qe*���
�]�;t��N�g3�Vg2;H�:R:邞M@��mB�B����g\w����<a����dӯ�)�)�SP�_2R��g�+�ӭ	<3��&k9�6`�
+N9>�\�lA�;���J�}��X� 	T�.R��D��@m�%9oFV�)�	��7���?*�
|� �d��RKcS�����q&�2�m:{7B(�RQpL�o�72Dn�^Rn�6H5����u55�m����8�}a��l*$�?�J��.�7`�$�4~Q������2�(4���Ē�l�]�E������(�(�������2Azw\�S1B�؎�����geD��������P#�Pe9Uv��	���e&O��H:�磲耿ޥ�����^u��A�G�{)<���M�C��n�H��rӗ9*�	$�p:A�4���zT���?��~�(4�.�3��E_���&8cgb���X7}�|���a�㥷Β,���E��сH����ohC�p�o��ȱ�cd��L�L<�t0@~���g#{q�t�ԥw'\e�ў��3!Qy�Ics�G�l��͊�@MBe韖̡G��\�j;��ZP�[J�JK+Ѭ�ބ�qے�8C@o����}����B""�~<':�1�.%eS�<n{r�r2��/���<��'�;�E�E�gI� �!{'��� `羦�����F�u�ծ�;�}'�܆J�BS�xϕA����5M�������/�;�i��~l�"�&R۠�X��wXR� T����2Mn4 ���h�K}4$x������r������Q}z�������c@�R���(�ؤ{�B�C|�7�_��s��ۄsͩ{��G�Q��<���$�E�L�raC��6g~��⁶���M��{l�j�+��]��\ͱ���<ŢW	�.��7aq�'�֦s�i���->�������q��}�|�TN�c!��e��Z�x�+O�����e ��[?����G���41�7sj�\v�B5�v#7)W�I�7
E=�&y�l�M�Ih��"OF��V1U8IfdaW"?����NL$�S��Ȑ�!&����vǤ��I/�`/��1����7����m�_��b6�>f��jj�0k�!m�����w�z�b��5�� t���H:�d�5�?"�� gZ̰iN���B*�>cs�:��o����c�eY3���4��xs{�}���kr� ���[�0��Ǩ?�������m�G$�E3���+�<?�������|�ٛ�ˬ��׭81��p������� �=Ws����o���R~��=,NKk�aH��1����~c�>�6����N<�Z���f�{��p��Ə�%D��K�4��"�Z^��Xְ#�W(�1�U�%kЮ ��>�c�3M@���J&���k[ڛ��5r�?��h�������m>i |܅y�zO���:q"A,�§$g��5̩ T.A��	x'�'�Q��9\��S�'�=!���e.�O�]k�����7��\�T�xf�+�$K_]�#���-zw��#��a8��:7E={"�.�q���1L̩���f���c�g����P�7zB!�f�Vq������ѻʴ��/{�ů���/�|���^��|P��R�Qo�4�!�ś�\�@�KR|�t4�_(]4�8Ym�W\,��3�fT	����/�Ԩ�%g{0��k��(�CS{-$��0�����.�T�`�;?7�>�U�f�U�6J�Z+:�C/���H�1"��I��ڲx��Ү"����m�� d�Gխ{*�5Ӆ�S�h�4��T�<Nhs��7p�}�d��H�Pb��a��������sUrLQ�h����ZR���7���ˬ�K�/q����0
�!�l��)��Vq�#!�	,7Vd�?$��������BA`��aF0)[`��n��oy���X���+7�8숶υ��p\O��SI���f0)>sw��{���10[=�n��u�f$�<1�v�*:��z��Ӝ��������4U�� H)��C��'��d��-7�뢸?��,t௣|o��}%�إ�~�^����|b�������s��$[[�J���v��,���=�_!e���v���$�X�J�)�����ScӇ#�?��oX�@[<4�����Y�?ՃU
�^��_���L0�JH��V\Y7b��h�"(���t�����@���聪����SFBr��,$E,� �[���������ae$:��e�>Ό�׵�����+�!�bқ�eq�=T�'�s{@��-N��kճT�T�d�����v��M��,�,�I��*�{"|����iڵQ况Ct3�5��	̎��x)�V,�� ��(�eB��k�G�^�}b�H���d��h��a�`��6�a�&=����<
`�٨kY��\�*[���D��[�|���p|�
Tm��-^��������t�M͢�76-�֥��"��� A
��l�$�S
��a���\����;�&�5�ͫ@&��ܘ=#�F{�r���3����t�@��Ub��Q,��4�y�M����B��w5C�\?�*Ϥ��Q�5b�`_$��L�I�G%�z[-.��US���n"vP`H��h{�o.C�Α��-�o��D=)⛯�S�
g
�b��8��\=��KS��
Jͣѹ�Yl&�ɦ�loԯ��86��ji�t�?�	�Ǚ�fl�5����y�+����M�O�%߈�I���Q�{�:��\gh#��r2X' ���ϵ�2�����/愇�o�L��հ�F�7u!?�-�`��af���{�,��0V݀�X���]zz�ɨ\@������	�c���C���	�t�����f��'>6GSM�
�ͫ�K� rs�[�߁Å<4<l��N�M%����7U�%cd��^�������X]h��0`�p�k�d't)����g��k��BA9�|=��/��}�2��7/tj�
rl7G,~����h]�|�8MzB�ԩ�i�T>���Ϸqaw�EZ���N�
�m𯰰WP��Y2h�C
�����>Xf%��%�J�w��S���[h�}W���=]`7��/�F�����hKNv��3T$'���#��9�Dc��!�U�)Q2�껝|����F͈�u oGk}���S�����O�~�m�O/��#�n�����G\�D�PW@k��u=/$�R�z���rP��-1��%�='�@��2�9W��G���.�zc�~�޾ym_�*�=����DQ�+'��22�EXg���KV4ˉ�l+C�Sń
�B�w��������=*6�,DS���S"���w���/��[,-��n}1��č���Q'�A�,� Z�-���:޹J����!��Bz�K�^�b�;H~�Ӷ���պ�2��9s����F��^��\-�o�
2�`UV`o?��S�@��M�u;ֹ�[2��y��f�3t�=�=H�22wB�;�I�kҎ	~����,�wJ"�'v�0 �̛=��5��[��	%Y�����������=d���
3x;4�+x�|W�����,"�٤���|ƅg�����L��o�C�{�5y�5+����5�?JЮ.7�t�3g�P���m�5��uD�T�Ĺ )a�M������XF?`���;7��Xx�ҫ!x��Q-Y�?;��e-C�	�b�٨�n9��W/�ѼX�A,tT	����<��
�1�Ͳ O^X�ik���y�.���R�BMZ&�=*!�R���9��h�ŕL������Q}�������yC�d4��"Kh�Z�Ϩ������i������U����gC1h��~i�`�%�N�4�>�¶ ��[�H�qIL&�_���:�
�^�o��x����}��$�o���QD��z�J�I]�j���$��47m�Pރ��=��i��:2����k`�D��N�!�&풀G�.I����V!3��̞}r>C7�}����K�Rm�z����{rc9���O��V5������iAã����A�v#V!zV���n���q긐��\u7AVqgi�!�sm�-��U�=A*?��u�����Ԟ��EƑ�z*rF�7|D�$pç�L���c)��@p��|��љ�U�-��e�y��J��R?��{�M���k5g�ɤlm������g���&�,2 z�o������,�ʩ��<�i"�A�v-I�ʹ���S�0��O���D�=^���Mt�i���s�2�z����l�z�T���9iQ����ۿ���X��2��e�=���5���=Y��IzU���-+)Po�S(߬����*����Q�;��J�