��/  �1%(�%º�6v&3q�[�bW�p8�a�7�Hԍ��g�B��J�fW�|���+S���EX#�;�sn\�q棘�-ܗ��i��� ٢z�����V�ZZ �0�k����S���ȳ�!�՗UM�����K���g�67%�r�E�EYu���ƥ�nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�nZ�iw��/��Ug����l�Ʉe����GzN�-�"��Cr����S,�d�+9߲��R�?I9Q����A��w5�����%���M�_.���)�`� �7C�/��Uݓ����i{��o@��RC����r�nm�X�q�1Ȩ���39���()���)"J�}G;� -�"�����	��š&�@L�2�E���n�kp�-�}��S4I8ı9�f-����4M�y���҅�4�JWw�g�"�^���v���v�i���A:���F`P�0�Q�+tF!��8E�V^{�P�u��_G��TrȷD�yO!�0]y�/�z��z�%��eO+a�9H�ϳ*�~.C���5�ֿB��ۄ�v;��ݚ���zUd%Q>����^I8Lס�6)#/���r�DU�'`�c�	�l��ػ+���{������P 3���i�w���*��� �Ը���\�Y�I���0��H)"�U,���Kˁ��mD@$p�(]��b�6%	�޵��*�?��2�y8�
�7�$.^P[�O������#ix�����X�3�����ҷ�W���D�NO���PX�U��#^Z;`���N5��=�DS�xL�����vj�I $����k2T0L�о�S����#���zDmU��������s�*Fj�&�GN~M�)��B�99�M���9��w��-�T�R��G#B���T��I#�߆ѐ~�_ tDN�W��v��X�0��R�ff�.`��m��2�ˡ[�T��8������1�CB���t?���|66Kr�oK����
���p���sF P���+�b��%��T��b�md)i������9�P(0Ec�$`zL�F�C��Q˒2�EڶI��_!l��_f�eҝ3+��2���AƤ�T���R�YPSV�����Eռ>E.��v��2��vӹ�h��es��	�#���}m	&$m9�ΰâx*��(�;�j����wx�q��\4��Y&g֌�7�}�e�;/e��w���7Q5E�(L#X{w<�χ��C�T~�o�l�s/� ���`�+qb��w����d��^�����`��&� ��;U��ɶ���/�I5���g��$�=c��R��ޝ�Ɂ�=��7P��ч�HmG�M\�9R�o\�Bq� ;�k�)��쇷����?��^n���7��i^ME�c����w�dK��@0<�n�kNy�Qwou�����1�.��i��)� Wݿ%"��=�K���v�}q2��q�?��X˕�?:r��"̻�w�+�Eq�;p&ڋ�V� ����qzL�*�B�=f�3��ͫ�Y��RFJ�P��d��O?Q��o�Uμ�(by�h�t$,�:\��b��ըz#CSFH� V6n☸�Z{b��\�B}N{�~�qdZ����Kqt{�3�|��^�?M��R��qѬS�d��+DD@\����\i�p�p� Se˥����4.�y��S�*��;$��Y8!��6Y8�������C���S�O1��`t��xN,�M��"M��k�<[&i2M��4{H��<?LX�rU��$"Ge����I.���qw-�i�z�Ci�ͬ��7���uZ(��V�~��i5�'O:e��dch�z�9ݮ�"} �n�LhJ���l�����giÎ��b[n��ڐ\ۻ�S�.tI����]���ηg�&mr#S`3l�~F<=����J�x���Nv�9�[9�!s�1[=U���蜊[	����һ��vXBڤo)ڡ̎��D��C��۠�8래��}]n���	L�X|t�f�z7���h��i�덨�8QS�߹	���S|�늺^^'����ɽkTr�.!{7�����Җi^W'X���&M`�6��zg"&,��~����w�����	�o��^�Pz��i1?��F��1��p��3���d&g�}���͓emW趣7���jmr�a<<3����9 � ��J�}���7�P�*S��=hȭ�C}�H�V��O�(�=m� �i� ��_��	@_ΰ,�_����W:e%6����ⱑ�������|���7Ja}YW|v�f��K��G+7`kav吮-�X0��{��u���d�;�K<�������������$d�t�-�S�g�R��+�����p�aAX逵K
|�9	�#^6�;䙑`B
��˪bE¾g��]��iS+nhL(Pz]P0���WO�Y�D����:������&50���;F	�9��k�������O��N�\Bh�8���x��r��rF9�}���҉f�/���B
��,؟��8&5�|�=q�?�����aH�_E��v�$���&$��E���w1B��]�������:�몷�E�C�z�Č̒V��׌��ɳ�'Wz�������˂+2- ��?W��$	ږ gFP�}�w�-<�3T��Ur� ǡ�� ������)�@P�2o�<F�u��f�җqz>���%�a#��o��sʭ�����>ҡи)n�L�Ԗ��MP �$p\ҥL����h�0ge�p=7�������P�cl�P�q�'h<�)Z�PW�L��q�U�d�t���X<�m4��3,��?M�����#�����O|)֤B��5G�lL��H� �����V^î��ո��7>�tF���-�pK�N�2�<*;_L3�+����(+���>"ur�b5��Lm���G�wf���V��jV˘�L����c���;1���t���&A���Ė����Q��R�b�����	���pj����knn?�Y��X&���,��o�����G!l�	�J�Q/�v3Ry���ߚ�.4���-�X/=jeG*,��WW������*ə5��r���E&��q]q=n�Fc:�ޖt�ċ��!v~�Ғ�2`_��i���k��ձ��g��$�D�|ȱ�ߚ�ރ�m�$���%��A����Rthƚ�Br��Hɓ|��	�v�%�ꄅwW�$�2�##NT2J��O��n����p�)1 ��s)0��2��2��RoX�g��2�o�~���r��e����p���#1O/���]9��A[����D��{5^/3�l#fE�wn2��ڑԣH��ݗ��Ng$�%Ǡ�3���A����!|��+�ګ2�V�z�?�¿�X�v)� �T�\n�=u)_̷�|��"�ET@��H�Nt�鬨%��'UP 1XBUCI�T09^�v���	�2�<r����3��䱠�f��vSy�k��M�QTϓ�*�<�d	�ض:���<Ch����U�(����Rf��\nP=�ϐ��	4/I�.Pݱ����1V�t��r\Ǳ�H�^���eKGQ�:��LOXA@��g���W�_��5Ž�=k4E����Z�S�@Æ��א�ʊ	�ˬ7�φ�IB`�겨���Wq%I�X���V�dPs��1�s�"*��#M�˖���r\��V��;ˢ���G
2W�/:U,�7�Up{�� "��D��;�b�}���w+�A���4s^�u�ش@4�C#Iv�$��n���C�� 7)Zaa�V��F�RL�������63���jo%14��}�P�^c�%�.��g�kcd-P�ݐ�J7{��X������ӭ:�%�87��4.�%Z��F����z�����^>U��*"�^���+�9�� �}M��]D\�L����(d޵���V\3��h��2Zy��c�o�����s	s��y��/��$-N��.���v ����A�{��U��2�P!Ē�x��z�n$�M���,Oϲe�0E9
��qu]��L����kgF�"=�w�� ez^��k|�Zh�⥶� ��ؕvv8�T�܎��Ɇ��yy� �[�	����\���7z��|��A����Ƽ"5#���D��)lgW�[R�uC�dXsVg���. �`�ʞ����� �c��2�m��u���~�s0�Ʌ���&Y��2o�1y��j��??�r,a���������r�05]�Z�K�;�ۃ*�<����Φ[�����!�k.%q�zf��߼��Si�Bx5BE�Y�0 �	���*;P� l�
q���Ԣ?�$1D�7U�<d6pI���g���0?�����PBw.Z魩J��3���m��(�g��ſ���.�A}�Y¨��J�� ��3�2�0	K�1u-��=�v̔u]3ǆ��-�1~�R_�Z�������./L�9ؑMmSS��;^�m��j
t���$?l����)G'n@*WZN�n*��N�*�H�txau �Z�1gO��z�OE4$���%�^�����ѯ���|BX��.d���g0�������j��]�������Fvg��J�zg�[�N����ur����h�L����HiVnʤzX��� L��Ct3g`�+L�����m�%��'СV���vE{�-�|����+H�}�F�-.��}�b����`ܢ$b�E�h�B��iWM`5��G�j�ۂq�p6�0�l�$�FBk�{�0�|�rɗ�@��������.�Z�O]��aj ���R�g��xS]�/�=
nWQI�D>���+��ЭT1M���ʿj@�l�`�Y ��ΎK���\��r��]�B����Kΰ*d�=Tz&�����o��[M�{
ꜱ>�������v?1��*2�e
F�a�jxR��h��%��XG0d�j�G����]�uO`Q�U������Hz�Rev�^0=��[n;y0�tڈЩLƘ��~�-��~�ۭw��yΙa�ze�2Ռ�o���:d�����k(�l��Ŏ� }#��ĕiV���l��B�a��7|�=�q�" �	ݕ�`r`%�E�>!׉��Q[4<���u�߆�_ٕ��Leu�,�>��<�j�b�[t���%�`���@$��F�R��P&��-�C��g�]V�˿�%��^�)�Ƀ! U����M����r{\�-��τa�H|�fh�Ӽ��.e����*�ᮓ5N'�6b�|-׍�9����Q�3@a5�Y��ES�W��<1���c���s���׻{-u��;���Zs��i��'2tCXJ�,+ E�:C}����H�QH�Y�@f7�b��r)!i���X���D��Ow���@]�:�|����L�փv�� }hp�>K�!�זc�؄�g���N�"��+�>�=���~^>���(.�y�3�1��1�~��_	���ose��_�s�5�>�YgJ��z'����L����j7��	K�F	�!䤆�C�P�T5� 
����Kԗ����o��RS �H���s�ᚹ�xj�����H),U7���O$*}E��!)�K���ǭ]]��H 3�tƓǒ��/v
�h�e�&��5��փ�����[Nݮi$��º0������|������-T5/���Fi�dɯb$�-�Ieġ/՛����QGFxL���s�ך��D7�S�<�9OR0Lqw������ɴ��);6�&l�}j���	6f>r1����0��|�ݣ,�pH�����F[ o�����݀L���Ah3�x�b�ݿ�R����u��d�Q�LCȓ��l��,噮�������͉V�Uܙ�+J3{2lE��$����u�|��*!d|+�(�0��3N�G�%'�@٣�yp�z�N:��5<����s[e��v7k�Hvp򘅲)��>@Ј�sL��C��7�i=$u&���5O�����Xm%��� BN6�7���Ԛ�Vܕ�)e�f���0�3�8h��H�������6>�٬y!�����e�T�v��p���Ĝ��w ��@K�{�D`0{�Ns!�e�b��������Q�<j@�	%-��V��nE9&*+v:���bBE�K�h~U��;�%%�~{J�r���
	�O�>K&� ��OB`�*��L�8��B�2���pi��O2(	ձܒ�=Q}<-�Ȯ��ݔ=�����O��#a'���"B'��f�m	
ܚU���7��� ��
V�'�a\h5���V����4��MC����U�HL�(u�>r��p���ti�&e�7�e�9嶐bV�.���aN6�n�{�VR�hzRx!�J����77I��I�� @�JOø�r��Dc6f�ڲ~��v��>|����S��2uQ���#�J�`���RR�_� ���AN�(�ߡ%"�Q�M�o(t	,����q�?'�,�L���l^h����{-�,xZ$�r]gg�&�
�20O兛鍔<$T��s�&�G�x�	��gӘ\� ���(\����%���`�dJjY<���p�⊁�D�Vrh]��thW����E
4�qk�ި"��w��xO�[3�fn�L���=�hv�m�)	�FzE������T-�q�:�&X�KR/-��S��a����l�u�N�����H�1�fuG �8�x�(s�#G,�MI_̻Nڸى�5��.ZH�&Kb�ຒm�V��@� /Qܳ��2�_0J���>�[⥦����4u0���+��� �k.���7]�yw	�����`�z"N���=�e˒6�}?a����XV�1�駫D{���I��Z�W����N��!�8`�l�����@$�k��?��L~;;�Dw<J1u�ɚB�Mv�Q�E~�)�N��0���q�7�ovи���肎�6f�f�Ұ�|1��	��6���łA��le��,�$�����r�f�bԡ�\"�H&96�[��V9��XV�G@��s��
��T�0�6���$�VWvX#78x3���5sgϊ5������Ho��T�Sce��_ǻ�qn�+3�5��+�{�Ҷ6P;ៈlX[��^3�
aN�x+U�"���%�̟%.��Z�����q{�!�t�BRo�PMُjvy���1�<�L�S�a1bd9����(�(��~�����~9��8�����Lo�ڣ)� �`UC���9�rI��z�𳠓��<.��K�%YB��8�x�\����`u��C�i�}�R�˄���q�i��Џ��Tt�������y,�o֮��#��b<�
�\e�*��@�f�I7-4�#�����s�V�� ϻ���bQ��=b,2QJ��I�c't��A�S�Zi�
���Ћux7���!?����*�A�Z��0c����A�/3 ��'�-:)0�#���U��z��.�<�:��`�S����׹�1��2#u��S,Je[;W�3t,��ί�|����]-\	�8/D�-]ͫ0��@F���~d���k�͗��SC����$�a;i�ǃ.U��WP
$�]�**`]�AM����@cnU��ae��)��Ӡ������~���`\�s	��F�_�����3����ij�O�<E���Qp
�B]�q��]�RCf��?�$�W�F`���Sk�i�e�aZL��T�J��H� {����x�\3�uR�'�i�}_V���.�"t�*�M�w�y�z��\^{~�6���c<oP"�?�!:��]��٪��Z6և%���X���ظ�I�\x�P	n�:1��=/��hD�u�`"u���¥;H�~M������W�X�rW�X��i�C���aZ 5���$��mJ!	l��y�d���8�r<]-�$_5���dc�F�dRvѦR6(�_	�� ��ކP���������	����R(*�XeD@@T�|�G3�'�G-^��v�-��Zp�°�J��m_���r��%%C]c�,�yu�Ϥ.����� ��f�)���蠇=�7X��PӜ����X���q\��*�Tm�ƅ�?~1����|�<(��±%�*�
9`|�EZ�Un�r�5Og�18_��z[���x)���K�6JL�E���!a���&�d�j�(^�{�D7�n��ۢ�1��&z	C��U�+yi���ąO����F�\K�^�۬�
r
A�aџ�xP�#��Ng�A�����k�A��������5���BӬ:_x��|Ca���~B�/�s�'F��2=H(s.�'�^vrr�p�dR�]F�������7��n�f��1����E;��_q]|u��4�ai���z��@.��=
�J��~�����@1��ֻx�		�`�ny*1�A�x���o�_�KtV�>���NT�� G8U��SIUz_b��b��z��`������̸}�਷9_7���~�6��a�	o�l���u���4��CE�18������;h�%c���P���],�bZ[�i��HG��ΊpK4�'/�ʴ�|�8�`u��P3����P�MVp�}�� Rn�ʥ�����E����_t���ۼ��%^��nm�unԃ���*�e>�_�� �fꀁ���4���70��LK�Ʈ\�'�҇:�c��@�y����bݹs��<��<��үgj��pI/c�^��푰�]7���DBw]��O��0�EE����l�n���m��2��:���`{7�Z��on/�َ�S9�M�	��)������A��̋.�/�j��~�}����A�@%�1�FC��Px&�j6��S�(�������Ie����<-��Q[R/��No��ex\f�:�i��G�V\��rZD��u����F�ݤ�� ?{M2��$H�Ё����Y���s���eJ]�E�a;��x�5�Aʇ��3:�����eweU���{�k�b�P��ѾJ�xY.�Eċ�*�fq�ȅ,���p�{-�!1	L>I���i��<�ߟNR�dyЫ�����M,a���1i�m%a�-L�W���y<�8If��e\���~�9t�uل\N��b�R�qx���0�
a�H��=��z��Jd��u�>n�gÒH3z�Mւ_1��UDj4��\�|㹋���W���<dR�����kӐ�1cs�u�W1g�&�`�:�a #������5�#�]v���g@�"�ALMM��I�s�zuR\�2_2�n���W�$��~�w�$�x�~W���D��)���(W�2gg1ռױ�7�1R��J>��L�����׫���UR��'1����wv��xk�
n���Oϓ��C����"��!2�S�u�*�T��Sh�i��f����sΖ��+aCC����:���qYCL��i|<^�F��I��IZ'o�a�(S�a�M����&�Рߢ�͕�S��O��Ѵ�[f�5	�����'�W#��bCc�$���	��o�w�\[A�f���[�yS@R���C��|zj��g�|���87���4�i�a��*��%Sx��?�4f����%�ӄ_E��'^�"N�[�'����)`��uY���+�ނw䰴�{��2�j��`ͻ�<�"*����?Lw���M����D�Ev�ω��aɢA}��L4t�~�g��cG �P��(������3� jD�fajzE��DA�cL	�)j��QP���tG��h���!��*��J���hCI�!��(�F ������S�oWZ�O`���*l����f��Զ��N�8�>��8}�UF��Ёp��5;)��o*�ݝX�SMn~F��S�3(j��H��n�p�m$W�c���1Z��S��=��y�$$/�Ѹ�ɮk���h�l��\XV�����Ǎ���k�����Fn��������:�'�[�:��s��ܞ��5�s��j�d�`y���(��l��xc�&�ނ������etf"�i���͓�#��6V2�����|	�p;���Ns��:Q�'�,(����O�7:�O�1�[m
шMw�@�iޡ��$Ί}1�j�I�6X�j ��'������ƾ��C�>�����R3�Wq	g�9�Ϛ�b�f�v���X�B��9<���	���2�em����j����,b��ó�a	ѩ���^7S���V��s���v��aZ�t5��e���� ֠��ql��e&k�f��nP�6���/]l�d�m��2��l,I��ep���-Se����W�\C��T�'�r�f��mҨ�t&8���g_�-�Zw��մ��߬\"�F�3g%��9�NDP��q�@�R��l�u����!��y�帓[
�k?1�Hn@#���u����Y���~E�#�4K�೦��n��U\ȮF��}+'<�:��oE�����x��Q�p��}0 �\�?���A9�iz����:)h�TG�Ot,�T�rʤ�\F;�|�yC�<��C��R����.�+�}?�B\)���y<��O��%J�� XK����f��ɜ%$��xr�O�\k
$�S���~�~98��,$�Ք�y�����t��t���hǕ��^j!�`����y\`̩�y�C���[t���=ʜ҆~�[�7���"���"FE�HM���}V>�j�4z���`mx!��WO�R�j�ʠ����ex� �������?����q��5d���s�ş��i|�)���V6�>OA�&@(�o�`���?1ؤ�|��_��t���W\ږѐOv!�w�v�\W�M�ɗF�ǰn���:!��We/���]-yPZP3'�;��0����>��.�9��<��?���YM_�)�!D���Ww��(�0q9Q�;um2��<��í$�m�]�WÜx���m�
���*3;?�����9�x�\<g�����9��۽�9�qx&N�W����)�>��2��9
� l�r��T�P��s�U7�V��D�w$�	a.M��5�JMgD��T�ZN��p��o�4��%0�*i)#�m��uHU˶>���o��:�ʏ� #�D����p�i��%gv�wjB�S̩�.��PO������^[$�P���F�|�F�p����'W?�"T;:L��B,Ga̵W�w@P-�>�Y�D}����#O���&�8D'�P�Haa�L���}�H!n�ˉݟፘ��"�R)��sq֌2�{q��u��Ȋmةh,�,{�f�̉����0J
��]|��p��W,;d�Ji��K�dQ��Tl<n�}�&;�)��ٝ'�u�B�п�r@8�X}z�&]JTf�����6�N`�T�� a��柈O<�/��͌������w�r��`+1��L�ķ�q9粇�������!R������0��h3*��ql$c�Բ�'&i�}�K[�i���\���T��az[$������Iw�]�gt"sK���/��X��%q��e�r8�����X���.{
��&GH��~�0֬o�Hz���Q��~��-�3��9���A��z ����3>�176�,���z�M�n��&F��k�S�B�ⵅ��Ϟ<ol��&��m^�"��we����2t�
r#�����+��t�c�'��B�Ai2q����f�P����x�_��!nf�>�3����g��K���	ىYr�,SAف�A���{`�� ��h-���$"$�>qu�>�?��ԶZPh/���Tw�Y_�Q����%س����*��a�����{����ʜ�h��̫o�1s
˰��.%V&����͟*�pR{����*�3��!�D���ƴ�8�� ��G�s�Y ��#�	Ǣ�) �0�6ЯE��ml���;�STB��/�6�'I�cm�Dڧ��K�y+iVЎ�s�!� ��t��򎐺�׺R�:�#�H0�d�jh��I�{B���:���O߲ʞ� ����`�b��дgH+��3p�]Ko��y+ ��8���iLj`��h��*����]�8I"I��/u3�H2���5������#��C�#���R9��į�sx*){�����T�!��,9iD��{^��퍿����T��x�9�RfjBN����Z�����/�l�]�x��\ ��?���fZ�����
�l�s�Ĺ]]83������*	�.2�Č��i�[X7�|1;��^�����A.���{�3L�p8@s�|���6?����R��,�
���<�u�;E��G�~,�N 
\�<�D�]�>K	����M�X@a�=��!�{�8�O��!�֓�7qڠs�'��^:i�<$���]���?*V�B����I�M�N����@Wyv£J���z�=���."��Z�a������ͥ}�{��$���U)H�x��~���3/>�zKTVr�JTR���u�g�����ң �'~����Ѐ��M�നn�41��*$���4�����9!��bfc4���U�G��YCao��f�?	��Ő&�{1�tB;���`�D�jŁ[�P�����Rݜ&�s)}��W� yr�L��Ɲ=Cd��^Z���~����Y�"���?j�ň�m�[�P��R쬳\�(���������v)�� �E�m���H�I༟|R���z2��AdoN�(M�68�G
����_K�ˍ�Z"�AgT��l;fkW�,r�����yY�	��1.W����^O����0S�<��D�&��V���3���d3Bf����ᛏ�_�Q+�K9Zk;��/�O��PWpֶ�\��_����<��a��P��o9(�э�%+ڭΆJ��3 ��C�+�
�G���aM2�Z�����?�~	nT�r��bx_�z���KAB�UK�zC��eI�ڄ���Ĵ0#�N*$uw�*3p�$����G�3�d��S��bH���T>�q"�X����-2�іU���@��;%����#��?���D暐��Lo��㒼�EU&�W枼���4���\q�Y�usJ/����ϊ��?�9Ӝ.�� ��`��@�\�̆U���`��D(b�fX�0�ڎiz�-/�T8������I��\�P򈽎A~}	N�����~��2QR��+R�<�P�ܸ0=�	�WUT����i��avd)>2�N3?4�'<FN���QV2[�
��(� ���w<�E����YmĹú:� ���l���l�+@�T�pws�����"�Ugp�̟�䊇?~����]�`L�^Hg�57K;�q�LV�� �7��A�]Á�(�i[&�kt$�\fƭ�D5CA��Z�ټ��e�H�r�w���o4bd�.&��ds�z��5 <��D��"N닳�4�gF8;��Q���w؜>(b�H�U�k��5WC������E����ъ�"�$NJ�dF�t��g9��BY I:>��q���~���pEY.�ݔ�bw(�Pdߺ��Gl?Z����)!�:ȡ��� �EhM~�3���^GB�6΂�{@��$蓸�`n�g�:�*��bw�V.�����������=�=��[O��z�M���g��`���o�w#S��I䌼
q�q�_�{�9o�b
�(���}����I{��+̐	�j��@�2'Y��ď�C�`���j�r�c�0�ܹ;�06>3i�RU�s�C��b(�~IUW����L�-1\a4�$�Ғ�Ṋ����[�P��*��g�ǖ���C�馔�)��
�C��TЏ��=i��B�8���@Jm\�'�k��k`�qS�2|�}D><x��~���]�#wӮ�Z���MG�m�[ߦ�����u��ۗ꺅��r'�$���[��x8dK�H�L���S˃�Ӥ��õZԅf��Si({t�lc#N��W9@�=�;M�䠓Lm�Ee�어�غ�%��p!AL��,�D=��0IR�v1_��6����}Lr{F��=(��ǫi�x9��{'L�����l	s���U�w�Y����T���a���6:��(�/KKmV���bqا:����5�3�f�.�t���0.�Chx`;�
4�����bf�qR��mP�q�Sel�G+�R��l� ���i13�c�376�y��)Q�����*���x?:����>�j������3�u�ͱ�(d��/g�!i����ĸ*+TH}ԫ���A�y�Gմ7����}�A{nl����Q�O���ɜ�a��;�o�ƥ_�*^ٴ�w�<X�R��7!k��,$��׮�I_�&}Z	�Ǭp���|�4%7*���h�����<�E����E��B��i�ѝ`赧^%ŵ�hf�[���� ĺ��5��s�N�}��,�$�V���;ǋ�� _�_�:�p�V
�IU��}���U$�Q<�(��U.��*�F1Ć����Eig�Kx�^���d����e�5e�|����� ��oCY�_I�q�"d� o�B�{�@�Q������t��+�KO�y"M���A�a�X���D�ژk{j-^��+mv[1��<�{|���ɐ$AcC�M���o�4(�4��U���,r��x�ߖMd/ �*�?J��(���ғ��b���4�to��XS~�L+Oz�M$"K�XK�,�-�{�6�2~S�d��;��� z����7��5�I�bԮ���ll쌓���G ���#Uc�g�Uc�^�.�XtX���_ɞh���uH�{G2$�l{&CC�O|��wh�-�����Dбm�B/	G�	z�/v��AF�_�f�8$��n��`�;�_	��"��	�5X�6��E��a�:�Դ���p���}�wr�p��b�o���uGOD��D�*g�\�P�z����R�=�װ7_�����Hʅ�.�[����[A��|�4�?h�w���"���6̮�"`�%+VcZ��.��qK�Q54r}���Q	��}n�#@�f���jY��^���f����\� ��d��-�73P�>�Kx����"�d����yd;��u}|�-�c!�J=�Q�S���Zt��O�T��F�3�����ū�1�=Z�K���N��@ݲ�A4�s�6�߾�<�p�%��ٌ}���9;�gp����}hL�j�z\���;Y�;�`�l������"���Ģ�!�*_Hh��8���HV�`����@^�%_�t$�IW�J&x_�3B�+�g΍�6�Y&/m��$�=�����Jн�aN^�m����IT\U���V �<��,�I��',m�l9d�8��� kBBΑ�P2_ ��ܰYi�u�r��(�0��-Y�/��+�r�Ա/�18�a��14xDAvw�q%fðL��$��֐�����x��t����
8k����0�f�jw�Vr�x���p@�U�\]�"A�k��$����}U�ԯ���]�͡;"Ы�bӴ���5�:�}�~�ڻ�~uj}�9����y?���18�kv�i^�����>d��<��sꫴ���	�����<�v1E�����m��c�o��/�z4*ne@r�'��,���d�j)r����J
EǶ|�P#�e�����,���;q��\>Њ7�VI�;V� �e�n|*�X(�.M���w�%�S�w��c9j�@���n���6�e�E��8&�֬��ⓞ�#��T�k#v����d��٬����J�uB�s���̯Q�N⹤�s :ᑳ3��Bp��%<u��'���L:0�.9$a�5�!K��z�xTi 2�b��`����X�����]h��pLfQ��������[�!��w9qطqyH<�o�3���f�0���ːЇ���64��%���lƶ@������;&��9Ӛ�z��"i8κ��8��tԜ��w���Ho��#�*Ϡa�*	���<D,�$��1}	ޤ��Ă�����������_�����+=2p؀��Y�I�.#y�;s��n[���	�m�7�8UX���oo�M�@�NOp�t{�%Z�X�C��[�����Ң�|�y3w�*+�o�a�#�Q�ܙ�ݪoz@:	e�����"�4
B�7��k>�7/��#�Og�v	���d;�]��e>�د��g�	WJ��I�����ya�� �P�� �@E44>��o�r>�P(�FB���<��N�5^9�k��3�������O&��A�ז��b�?��ύ��������v�۷+у�ݜhL���^�>�_sH-�!�ׅ-��^�nQ��d�}	9=��f��RKf*fD\�4�ο�T�%�$fI�R,�)nC� � �UX���	�1��|���c�h�:�z
=G���	���u�
�"Rx��48�.e~��DyZ2��3�{_P`+y}5����qL���u�����%��a�!�M���<��0����=�����&�7��j7"�:  �O9����v˦�{ �N�p����f�r.Ѕ��g�q�f�_ܢf��˻D�6�����5}J���I=�4�a|����1�ʊ8.�g!�!�e�[W�����,ޛ��l�\z�t~cCLG�ž�d�0�j@����Ŏ�.��9���0pi-%6��:���R��8뙧�QKЩ��J�����:S
v�SyAaJ]�'_'�<���ŀWo0���;�q�p�*��4=�?bU���=S)k�
��k�V�
G�,b>� �ٕ��b|��I�X4�&=��9�L;�w}
~���4�
F�o~J���yDu�B}���q̄���;^A��La��-��$��D���n�X)c����P�Zy�}�?���a�Sy�*��-��GZ��Ҕ����ֳf�$,�M�ؼ̯R�T!D�wʮR��SM��b���)��i�w���@r :S,��Td��m��>��l���ig��ךm=�p{·��+�w���(7Yl��"eWk�$ �c�z(��^�������e�� �XЬx���Ѝ9��ǖ�Dpf��Z�RK��֒�i*0K��L]��h�S����H{�ر��Ynq`/R�ح�Y�6�6[���RP:.3��jtx�������|��+w|���#�Om4[�>�Z�W5��x�r�SL�V�w%"0��E0�[J6!!��Y<�y��g����9%�E���J;��������Ly>��]�n�$��Ϊ�Wm��[��s���ו� ��*��<}N/�]1��Do�PQE��G��#��{������I�t~2��~��x,5jQ�w~o&)ઙ�g"K���7��S��Oc�\y�8��{��?V�
�D��|["
�c�2��4��ɵp[���Ma��/��t2��!MB9��Y��ߏ���v����U�x�L�2�N6��\"���G����Z3�9���mw�B��FJ�8��Y_(���a�p�((���<~)%f�cLZ��~�M�9t�]�t5����d����oe�H둦��Q��оD�P(�o�ד��=�	]���!�aU[�"{'�?�c�
�6��F�7?���0�~����! �*�������iܜ^θ8�0RZ�4��׬i�6}9�d�i�U� �0����8ܽ��p�݃dф������{!�X50�]��T�$(A����<"
�mz��4d�����3�m���w)ڗ�a�x�Oe�7t���]�"S,/+�m��"��N�}��G�fG^I���!wh�5R��Z�fO�>�$���%�����O%3&�HWЧ�1��@oy��N��u����I����>eX��]]V��$�|��9-�Bk�E�}�y��OY���%�`��V��|�l�"H���$��p�M�|��B�_��~b"��C�,l�fu�U��.�{�C(���-ɴ��!��qJ���d�ܝ?��Gk&��i	"cT�]�Wg@VR�A��&�6>�a�%�j
��f1�������#;���",e͛��Xśϐ�!?1��h����,��O�@(F����X�H0�]�}�H5�+�P(�TD��Oi"|.�Ǯ��6������n�B���pg�Vw��*������wC\�ȭ�R֘f�"rvʜ#�8S�[��]���<B�;0g��9����D�ѱ#���7��+M�'=@c�*�W�)�dk`m� d�M�&J�/�m������=*-M$^��A��I�hF�	7}-�����V߅���DKV&O�D��z�l)h�����%���+��m�V��C�����G����UG�>�2��Jv�����,[�ʷ�"�f�+?��诅�q~�{{7��{�t�^�~#�~y�C�ȭ�\8zz�g��)�4����W�s�}��'����j��&ʓ��2��o��[�⧨�E��7?D>'-�T����f��9+�'�"h��M��C�����.�R��AZ#�'>��c���tx�B6���Ziܕ�!��
�ݧ0_���`�7F�Y ç�$t�+	ݴ����p�g�9�v8��y~��LA�����t�R]�ԙ��3�w���Ŕ��NOTA X^'V%t]Hf� Eu����e#i�����qw�C��������#]PV�����˪3�\��ۀ<��M�}�p�~� >���f�Ui���s3e��]2	|�+�"[_3�J���n8�orh����[��E���M�%���g6��i-���9zm����m1M�r�9Ԣ�xR���_����j�h'9��YԿR�l��������&�#���9X��yf�n���п�R�g�Y�$��ʰ̎�gر�6�˓�MS�\��_+���<��w�"��H��rG��t�7Eb,�fX>!f�"������(M���Q��Hu�L���](��~����Dr�|m��A�L�U�!)^�a�y����yA�5D�|.)ejx�w�qG[e��i� �=k�5=h�>X��5���G=�{��t�s|J1I���gEs�VCȊvO��!
ǏƆ�I��8���\	Y|�+>2*�{E�JyD�E�w\*��N���q��]q	�X�^Hi4�
I���zh��;�ը:�q��*%$�U�Y�G⩇7�RFZ`r�y���t�χ�`0���1j�<�5��0��sZ8f1!jٵ����yq���	�|��e�k� �v�o��H �������\�}%��}�a�O��lG��|5�U��?ҰKι��+�q�%;��OjCs�*J˪��/.��٣���+�E,�8��H"�(�Y�|S-��V��g������[�cF�Ѡ�α�5�(�j��ҡ�4͚%wr�F��1����4��m���6H���H�f�g����8V�v�E��-R��GZ��=��������33�9�2e�/䱅�Eo���dQ��=!��A;;�'Kp>Y(��w�I>D���f.�7z���l:@^��8�^U~���hV�%�.�|�����cTEU`K�w�X�'v�[�#;S!������mV��	� +���%�(:��p:�p��S��\��d��lݵ� 2e7�(pm���,�8Jе��̃�_�a��-o߇�X#.fq-�l&����@ᮔᅆo29]/��jh�:�����a/U�'cXQ��2�2r>R:�K�8�Z�f �L�; �q}�G�s�F�X��S��Ե9��+���}d�J���_��(8'���T_v��?�"�2R��!XG�g��K7z��}~\��j�a���F9mx�����˘	zK�"d��!�:�c� �pA.��qD:��&�ȒrbQM��]�ӿb�*�;�C�,)�q�/�R�� X�S��W%�W�Ƅ��F&:
�h�_`�f�qF�O����w���s~*�w�c�D����ADWα��|f������5֐%`:�!��L������I��h,��C�ѧ�*�>V��_�+I6?y�ߨr�y��}�����5P���q��罤���czW_倱MצT,f�RJ:�v�A�x Ε�]�i��Tr3%�� ?q���'Ql(+#��r�A�Z�y��n?q�6ѡ������<�OX������QI��b�/rHL��H��;�Bc̬�z@:�مE���6CGa2�����?2)l���p5���ܿ_��0� �V�����Fɍ4��.�S⵱��,qv�Kѭw,18�xg���'�B�MC��N�5��\+L��R x�=U%~�z�9����v�Rѳ�Qc
��������ӣ�]+�26(�B��6�������+����k�tY)���G�����hX���o�	>꿫��(7X���=`���s��4���C�ڗI(7���A�����H�`��m}F����#��1��1J���+.	�5;c41�kY�bf��l ��UDy�p��#�t�"�t��3�J����Eq�A�F��^]��������p0�k#��:�ϭѹf��a���RG��ȵ;�끋:v�3�1�"����}1�{%�ƣ+͵��J���E�f��T���T�S60�X���u#��=��#��f�$��)Y��}���G�`�6����8�o�S��	
�l������7JX쒖3�0�q=M����N4޻���;������X�']5#�1S*?]�Gr��=��
�����-
N��1R��-��"�|Ԫ��x�q��
+&3���B©mD��ř��#0�����j�Ѣ��w��Iz�"�X�y�9u�+�2{�Xᆦ\�:���b�wѾ�YAJ����؃ШD�P���<�#J�VQ�a�}��1���w��e�`I������:ͤ.w��#VaZx�<��nG|���sv��%P���њ�ut>\��ө�L}Q`��"�x�AZ�~~�D��#�C�sN��W�����$�6+:�&jy��	r(p�����:� �Q�3� ���W���B��>_�5ʛ8���7��֏���-&�Lh��G��ֱ��V3�hgm�\S,�N'���n�|B(t_e@$7鳭9]��-�1 � ,�]��Ïh1� ���(����n���:ߕ}W�N�h�[F]�Vt����7�	�H��l����|�Ib6k���M��&�<�������c���ҵf��$�E�&�����\�s�ߤ�f��@b'Jd�������v��0��%�Oi<��&���P�������O�4�ʪ!�N;���E}�cL�PW�SkH_�)R$zAo�h�SQ��Y<��	8�ß6
��������M��M�@�p���^$+�B߷�|ԶP�c�32�om���-rk����+�ĭv��EO�AGu`P��6j�n�ӍI$���F7JIǖR�u�qn��<�!1y��뛟�A��KO�:�_���o�a"tc�F)�k��C��I �K�9����Y��0J�����B�g]Ħ�������e�+?v=>�I�Z�����!;�����3,�t�~ 1�*T�M}+����w����>���+��Q�3GP�6�Aɕ�鮇�~�q�Q�0��Koݰ-
q���)��������Z_����5/.��+���M�fپ[0�F˒��H�1>Y�ty���T=�:zK��7"��	���N㪞UM��8l�z��d(�/Ƿ���w/�TZ/�R\;6�@�gl���7�x��c���)�5��ڻj���8=�X9z���s�8�K�ʊ���E���ǭ���M�	p����wa�Z��b�
�u3���Дʆ��nm=AK�3Z]�a��I����t�P±?
h�����b�U{��C�7���{�ų[$�I�HX�7��{Z� 7�禅^Xj^�v��x�%�(t�;^��Ҋ$���˪��՘���u���aB�C�i�qX���s~J�mQ�G�$�S*Kd�ߋ7��.����k���֩�l�G%nFt�p��������^ZK��5¾t��W�k?øI�&�YS8���T_�6$��f/j��F("XBۍA�h��e+�{P�����[�-^�.�'�x�h�VE���&�h��;����������A�셒����������'4�����PE�륮�a�Oj�v�b�R����jΙ�6^�����CdX���3!��b��N}ń<_R�e>*{���Q��Gg��M�٩��V0���|k��~	ī������r=�����B.I����F�FvӪ��Fw�Hq�vӳxhlψ���{N�W0���T�d�Z�Z�M��s���G��0gr��i�H�������n �h�h��_��ML+g v�c�ݥ�����jTΞ5n*�}�(&(�/���4_�Pw��	bj�9>��&dI=x�+=��¹71@�[�'Qb����0�B��قnL���okV�"d7aD�vAe�m��GL('��WY��tݒ[u�Д��yG�m{I�PQ�]w��'t@M8j^s�m�ߕ��EЯ��U���PG��]]%�.�6�}�$�K��S{ɦ_��[#��X8qsy���A�t@��'����ք���$��E�~9��~
�.�J~dV'��Ê����٫�4W琄�����4F=����D`�;"$�|�K��և|4����@&��#�D'�vj��]�J��r#W	d���k;$QQ���h��-q���J��ܘ��hn�.3���a@}#.XՅ'C�e�Д�1<�dc����1�O*�i�C?ճ���Q�\����l��)�i��������Z#x�N��-��A�#���U6�j3�˚�����ii��s��J�����+�w�uF�*�=�L	V�;�{��w������cHe@��}+�n�?�H�V�5+��J�Q�A�>�K-�a䚖vH�I��nd��P1~��1_»cwL�Z�Me����>!�;���� sOZ�����@�Ϋ�N��h�"h�D�9�s>�DS�[5ԧ�~�����q��k����ٔ�4���f*�a�h��*�RP.`s��3�����X�r7<Ʀ3bj��ˑF����@xQ�A�p����-������$�N��гn�(���rp\��MS�_O-����r���c?�Ccy�B�il�j��`
g��I<.� 5_N�L|FZ�m�f!�ѹ��Y\TN�t�p��D���Ə�I��02 �5��l�fK$�aC�ig7�c),��Zx]��E7&�a_�tsFi/±寊V�1�f'r��f��Ⱞ����ۅBˑ��m�[�n^���(�e�����t����y��x�:��2��E����p�wKq�ʡ�u�7j�0g+�(�B�����e��d��L��#��W3�)�7�t$GP��d�q$�S��fF�����w-vF��
x=��3�b_�v�cA�G��K�ᇼw1��٤&7���_(<~B>]�k�czja�VXqԤ���]�<rlJT�<x��2�(o`	���L
�N���!]k|�Jn	���T)���?�@��*�}��ƚC�^B�.Y��F�k�;q���wTX�߯�j"[n��'�'�m��Ĳ\�I����w@G��V�.H8ʵ\r����c��u�����<���*�6���nA� ���U�\��>E�s [otΦ�SLl�sD"���X��l�C�������zoυ����@(p�Bξ����۔����J��L���X��|1 VF�<,a����?��7?xVItׂ��P�ՙ]R�`қ%���q��Zw�Q_�Aéu��?�h���ו}!����'�6�Y��G�nA}�{��ԙ���1zܡ�7�I��'w$���#`$X����V�C�&Ի�Ì�HdSٸy��^ǯ<%�r5W�#n�y'��h���1)���v}+:ܣ)�n]�S.�.d��Wc!^!Bw$R����`�_�.e���u���oc���^4���e��d���mW:�f�^sM9�I/��dK�hኅW��5�������pKR����ɓ��6�0c�`�8r!���2^�m����|�S����D�0��o�MN�q��Z���C��'�V�����w�Z	�;�<�m�q05�D�2��>���dҳQ�ċ��� S=~�KGi��Ť��PZ��fav�b�p��c6�dm���R�Ч~z�w��rֳM�(1�iǻƺ~yRS����E��C�`ݣJ6Us�/�#���$��{�0�����t{��
[!���1�}����U��>��@䟀�����e"�nQ���C\��A��E���?�k;�v;��Vڲ4Q~ļŹ��Wo.�����/E��KB�Y�DV���9s����Ӫ*ɰ5V�x�R�Ff�#[�tmYd۾�_��g�V�.T�'w]��R6R���n��V^���S�?갩XV�SB	�/)Oؑ��H��C�t��Ki<e8W���%���H�m���̱χř�%��Vd�<��"���������rݬ��S�7rR����6H<�_(w���&U6��S���x��ݗ\Pg������y��]5%6J�"a�{�-�঩����yX��ԓ���}9���ٱ~��./3"��H:�h�f��d�4v�'��{%�����l2߼�V���g�?׮�QP��/��l��:�����"S�b�����W�j�13����f�y-���dH�W�;2��-�ñو��΂����g���۵%�|2���ax#�`]c�K��[�,�!g^XH�+���:)5��ONIb�VrN�s�g'�
/6���%ק�7��,�L����:zP��F��L��p��l���Q����O�2�QB�0Z_`�A�lz>{*F{)0��Ey�ל�~�eT���/M8 c������K�k;���(�?*��)�CP
g���ڹ��W�E{�?3S��󇫠o+p��d
BKx���JC�Jv���"�㢵>�B9}8L
<R:V��8�ˠ"�j�g���I�7�R4r1�Qd`��]<zެ���o9�QZaG����[M2�QD���
�)��>��IVTY�b�>y4�$ֵ�
��L�(��~q�Gm�`���F!޶@m��Z��HK�cM�\z�VCej�?E�e��E/G����_�R���j�����h�Dl��(�+ޙd1j8e�b��.�y�Q�*����9����=8�~K`3�dPj���Pۄ���+���yʁ�/ ���yM*�}�p�������tڒmQ�R�#��Oj��PL�Xv�����L���HQ��>n	 �'���yU]kꍤ�&wA�*O��J%`�4�A7ujB	F�˹�ɞ����a���$�>`Zh���©�m�~��[u��N��P�1�?g��e��Y���8�"��1}��)�.�Ǻqo`�p����ɪ-���}Y��徜��b�	�\m�k8'�Ebw;|�c����wP��fw�Y��{�LI;�d�؞P� ��:}����Y�t���<k#�8�{ja!��?+��Ρ��.�8�4b1(�59�Xx��
p�>m�Z���w������)cw�ס�'�����;��p�& l����}�R�f`�]�ʃ�鑈��AO6�liB�/��h �U���(Vz�ӟZ�n�@�@ztȮ�lO��Zp�5�#Z����BӦ�4i� �����u�+l]M��|���pbۂ�M���]�ǉo��a�9R���=�A���G�{К[&0�1.�q��������d}�aĦ[��eAn�e�6���H��v8�\��M�eU�X����eQ8�C2��*�ޅ!�4���ȑ�G�Y��"XY�b%��tV@�n��Ӵ����
��_�����(:Lۇ�S��Q4U�X��=]�����'hZz�i߸豊䭍�a������0�����rk�����S#9]{d�eYP��|4���0>d,Φ+[�]ۿO�!�ͼչ�{�7�(f���"������w%�%l���A���g)۫\�8iVP����EC�{ϝm ۗ=;����yf-G��s����n��0�<f���]Ma�5j�q��㲻������c��Y��K55��޽�s,�r��;w�
"A���+�"�< F�M�AU�lL��m~�-�l��>�D��;�T�E�?�_o��?��π���u��2Z�?5)F�����Y�3�ꐔM����54wUj���b<l���;�������Z��/E�[Pg��"n!�/=����w�{��x���m_}5���l���
�T�.;o�qT�t�=������<m����!-r�[��n�h&�jw�� 6���Q�����CD7��Q�͹��;�z(qAD�86�8�Ix
׬ŉv�;ɵ�T��jA3�����XS�L�K[ d��L�+�r�����L��`{n%�9��z�q���V�s�#e��W�Vm`{���0D`���U�2ĥu?���&nw���\���� ����P�V�V�q �h!�S'���aMLj��ث����	A�`�%yd:�X;���JO=2��8�,�9/*715������=Y_}���9}!��$�̻6���Qw�L,�� J~��ϥ�&���켋(��p��p�%�|p��r4�jZ�M����3 Je��K��%j��Zժ4`/n8A�q�y4�,��Փ�B�8�(3NWۧ��ʒ�Ցgt�������y�TY�ď:���~F���2Qr*�o��s,	�yJy��7�BS>�P'��5�b��tG�H3�%7���-���������E��0��0�ʨ�.���,���Q�X��UC7�@`��r�T���n��SØ|U����n5A��p��L=�~�_�e"�>�E◷��6>>�	��tȺf���l��z��*�^o<1�g�b����!��QX8Ǩ�( ��G���M���e	���\��?L)h�?��)���$��Y��&q�Hh͔��rd���.t�H#��G�? ��iA����S��eG�*���%��m��q���u_<Y)=xz��m|���-I�+"6oD��V=Hh�u?���h�j���ق��txo�l =�:�d���w�M/�����m�A˖���.�ؕ��E����Ul���>��U�F�O=���q��J<CD��srE�	mK�����5�"��X��/�������)$= ��I�H�����%L�dp���M�hJ5?�4$`@�z�j�����,��v�p���or5p�����~�%����R�?5!��ު٬#��c[NP�L��\Kt�$~V�ޥ�
$��M�X�O�
;�v���N����+�ǳ�sE�� Z_{��:��U��d�ņ�����ԏtX5	#� �����A��e�����P�@HP( �x�¶h��s�Z������Ss
ŧ�Ē��AH�����ȅ�Ѓ���5s>8���c(�"�P�4�4��G�/��z�U��(�����n���7���c���wG�����n���(�q�I�dD�
N;��e�G�QD�Kv�V�ێ�
�w�v���k�@3MjJ2Zg�b*��ʮ]'+	v�����
�Z� ��If~��-N�J9�7����.4��8T�v���T��2C�2`�l��n"&�����K��:l��B���$r�J�.k���7�+�k0���
���y�J�T�[e��Bƥl*G�}��ۑ�)�ѓ<ay.��?C�r�ޞ��A����2&R<��N��e�r	 78BW���Φ�,돞���>�e�q�|�*l0i�o��N�Xt}����у�Y�3�3�p�-GG�e1306A�V���k`�`�8�)>X�؍�,�]�dzkY�q�����DX5��1���t����ݥl�0����`߃�W���N!o���P2����1l�N4��>�Lw������[�H ��݋w�Z}���^s�FՕ�	ɢ���'T�kL��@�B�a����9���Iv4]X��%���l�޳^&a�#͗x�S�GO���馑r���,�X5���⮧<��t!�j*w��X�;��$�F���\�[֐Y�o4�[4�D13�I�)nz�巭92�X |"�r%z�DU�a&��c!����'��1i�H2Sc ����eW��.���b�8�3�+�'Ŧ�x��镊�v+v-szq�â�>=&�{<K�=su��ł��w����iJ�cl�d.[�N�X����(���d�g �&�?�0�i�d�Y��1	�p0J0\�u�8�\W�<o���.�un�z�bc�+&��l��m|	����w)�Y�P?*�ZH���O� kUw��T�y