��/  τ0(]Tې��`l�j����Ry�������7Jj}�O]������6�i�<<��i�e��	��탸�hs�����-�v��	���;]�0U�(���~ZF����)����t/����q��mV-�u �z�����[�u���0͠��G*��F��=�`����nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�nG�v4�iZ���ÔgVwC/�N�T�_�;B���vQ����B�J���/�~�V�Iڪg���/&c37"+x׳�G���E����<�q� �^E�0���YA�$�� �U��BAp��7K�.Df��D��X�܌v���(����/Q�a]33\Ѫ3�t�5U����|nVm����t�e#���f����Q�*��WP^���;��M�m% ?Z���(�CO��k���A��G���'-���H �9|����N�������L~�/�N���p��O3��VU��Rz1X��9�W�W=k�[sre+p����K}�P�g��ow��#��*"1�D���4'��j��%��a�GD�m��ڭ���M����s�K(����^F,}�.F��3����W-k[�ٓ�!k�R���p�m0f>;�]�dʞ��jo~�S~��\��I�����0&�=]0�uU�i��GF��%�vu�X��RHgX^ܿq�>��6.&z<�|1�����W�u�YH8ӂ�rp��
	W�q�zU*�U��xk��ڥ��7U����=r��F�8�������[���8���Ѝ�uOOW��P�^�6i���+W�m�WgZ� d4��p�ҵSJ��ƪ�kg�&�c�5b��E��w+T	ꅛ#��f��%V�dC��_X*b����%[#?��m���ܘTr:�r���e��z5#�ST�d���WAz{�2���؞��l�%P��Pf��^~�ټ��.SF\��D,@|��x#暈x���.ǋ�Q������Q�������I����[&�I���0�NT4a�O�6�	�{�B*L�;Ťۯ����2�m>�{HR���s�R'�U;�Sa�[p��F�}�37,uX���<�:�fO*ԭ�{Ra�^{�#6K�K9����MO:�^iʶ�q����L)r@X	o��lNnN�ցɊg��u�=<y��g>d�# ��^�ws;�0�u;��Jj5���p9��y0n�>@̜f�1�Z�R�<	�g��.���@Up��(-tH%�#�8��dZM�Pz��׷Y���
�?�	�ov J�Z�*�@�D�窇�=f��c�d�B:�Y�pD9�VR�����{�"f��a�(�}L�0��!�B?��
���%L����w/���e�-�dD5���i̖?�L� ���.3K�jq\�*�j����)��M��y�Q��D نD��u;0F{�,'����{��,FaN�Uc�z����{A��{
�T��M�F����׼F�x,����j����j9�������1��
l��4���Q�)��������x��*?�W�9*dU$�X�BYr �y��"��2/;�"�"��{j�Υ$#�������V=�TؤG����Ѳx�
���K���Nz~.��-P��sn��>j7�f���)C��qf��~��r�~N	<"G-K�c� 2��x�9��҇�[ ��<��驱��<Sd�>��ubW	���_DI��s|=�1�rf��c�w6�_��>R��3k������T��U�0�=س����ISD��uLFN!%���r���+���F(wґ�9�_ H<�NS9ٮJ&���1󄗾>za���|��c�G�[� ��>y1�"���{o�?��]m�V�#�����x��0�����n�|���'}V?^�g��%ip[:�,X=�E�o ���	W��-����
�Kb?�)��Rh�F��I��ݑ�*Qw -�X�x�Ǆµ�A��-��\tw�r�����dW�`U���F+�c�#��۫�Dn�����Θ��wZ�S$��l�eu�R�Xj�[A�Rylx�u&t!�\��lG/*���p��9<�/{̎�mi/�3x(���t䏖��12+H���SӻtI�x.j�6W���jW���̏��B��Ә�4��9.=�\x����N�h^y<<�9���I�"<9��",���r�R�k
�?B�^���U��sQk;nO!���p�pd�}]�M����o*O��$��L[\�T3��qe�﯑�t?P���
"��mJl��i�/�]�1�B��y�,��tnev�V.��fX}`Y�x�����Ao��u���V�||p�o<_����������$��ͨ��BNWLQ`˩�uUR�ml1��NΎ���5��P×o�_kV[jo��'4io�m~k��L:ݏ�)���4���>C�Ɲ8G�6J�I�Jh�:��:�mȩ'���c�V�vy��]�n�m�SW��O�lq*t;"�X+�y��q����oe�*�$��WQl��D�4�,����J� ~�mX&�N�1K��\J�L��V���(ż�[]!���YK
��NeK�$G���+�`1��/���F�~^� �h�t.�PN�#�"��)����BZ��x������ /���[��c� �W�@�6�k��}�Y\Z<b����l�ei���~��#gឈ�?�Ow짮C��FT��f#;N��⽘�A$���W��ɏ��v~G�-�!l���mW�dY�*�H�v�yQ�a�=
�H�?�4}�n%	M��+�К}0��ž:�ʦ��k��]|�X�z�X�1����<����/�\z��6x��tt��LN����CT�ETT��;(
�7
�0F]��W`RC�F*�N;)$�y�z�$�r�Aa<^�4��><���p>�1��"<z�y��Ƀ�/���8,��؜�e{-V��NՍ�+z���)�i��6�P�"tv*��~y�Xk�����΁c�.,)��:��XhJ՞����B��4p��8�E5��1�.$���L�<6Q��\�&xt.hdnm%�)O'˻���������:�,R��^R�O�t���B�$V�
�iSc�xty��mR�@�
�$���, 8�[j�A���`����9���ܱ"�Z|`�$
	K��)bOhCi��T��A��NS�5��fe�Nb(P�ؠ]6�]�3:�^ٖ2t�奭���B|\��8��+��\�T��pm����(��u?�=��ȫC��Vx%3밚p�o���c����������ua|����|�m?&;4�N���8���̕D^NDZ�7&wUL�R�_�N)7�m;�����<g=�M���$�LN��W�T�Q�E����u}��
��~:�蒐�@�"[�~���)GA�lxih*�I|�w�R����s�m�� �Fڟ)d �������X�+��}D�-�lO�X+C&	�T��[D���H�5Wx<��D�fLk��]Ck7ȶ�mQ�ۂ�E����B/̦��)]#M�Nck��^�N�$�@ʹ�+��	���IK"�NQ���=^����T_����W�nDOJ�q���jx�V��
�Zl�L��\������L/p�� �&^�2�
����f?�7����n%_lO�4C�������5��=���{ȱ��<�4�����B�D����mƱ&Dp����Oѫ^��7�1,��f~���$4(�U7>m�)��u�w�07{YT�Ǎ�*�"C��9@���-z�#�YRl��%ʔ�h#N�j�

-���y�5O,v�6�,$�@Q�t��u/|t�D�g4C��Ԥfą�A�(#h]Ue�惃֟h��&;)�!n����+4 ��i�L�N��]�7z��������b`��w��z�����<Ա�h=�$��ڙ.O����b�^�����2໰" ��z������;�����NB�i$�A�7���(ng
����+b��Id�	��x0r#�����g�3Li�f���}R��*h?T:�ڈ��ɟ��!�^Њ�O'�v�r�{)�s��{c��6��ݨ����s��ۉ��B�c(M���������������7�
Ï�ۊ��è�y�h1����h����p!�2�9�h��@�y�qD0]Zb;�C�!�mR[j��m�.�Dq��
bQ�v�-��SJ���
R6+��좗�.{��}wi�#���AE� |A������[�Go��F�g�P=6X���%�تE�����Dy��nmZ��6T�'���A�UJ8��8:�	���Q�ܕ�ĉ!m�4g���gZ��m��Z�6M-/�#�����r͂�8�;2������v L
�0ݝ�,�Y#9m