��/  �^���H����^6o����F���k�5��n!ͱ�.䲴�w^ݲ��Vk��XϏ�P9{)�l�ll��oDG�Esx��b+����>ܯ�(��X>L�a%	R�iFO.3ѽ�sa��˸+���6qsB��]_��
J�W6��~*`.$�{�z���B%d�Q��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�nG�v4�iZ���ÔgVwC/�N�T�_�;B���vQ����B�J���/�~�V�Iڪg���/&�r�r��I����?!�Zb��{ �B��g�Ov�ϐ9HP��@�q���)��D��ͫ���t�>ND�[
��`	�x�Li}3�Л���=`�j�����'|��Q�`�f!�%���oҐAYWe+]ԓD��۹ڪNjT�Wb�y���NN���N��6�5�lI�aK:�Dqn��v�/O/�I���J�.)�a�>�O]"�8�H�E'~L�ؔ���w���W��M��-���&��虊��D�͈Ne��K�ڋ��Kw��ʾ�xW��-	��N8ލ�s��̝~7�-"��ד�RM��yK{Ag���S��DTFE�2�Yw��x�{�����?<{�Z�fvFae%�j|���h���I3���hGq͂3�(Ծ�ҩ�14�u|U͝�/T�;>�gL�a���-�BUk��,\�0Q�����ժ|j���dvS5��3��1�o	�Bk�Y���]Cgג��k�?��H�Z*RZ��:¸�?�p���3��C0�$)~�X)�V�E	���ʴ��ї�_y ��{���w�-�%�P 7rh�'�}�ySR�!z_J�(k��lV���w�כ�W&R��q����]��� v�c��3GɄRY���h�&((�}�'���1awg�:����@�g,���axi7 Bs�¹�sm"J#i��ū�Q���Ʊ��Y���,#�v�ܻ�Xe�B,4F���4�`ꫯ�t�4��Q;�s�,��$���ce	XyY��JSC&ʩxX� ���� ��m�_N��s�"-͹uu`�=��'�(�0],����[P;3�%_$w
}3�V��4�U�SםL�CJ����K����f4'�MR尅JC�F.T��x���Rw[����>�v��Wy{��yÿ����X����B$jʂ����#*��Bl&ɂb`��\���턂s���7Xc����i+�ښ�rC\�SA�>�Ф�bI�T���ME9j��FoQ��&ӡ�=�Z�7Z �+[�G|�5m�����y���2t���0����my!��%Nk��#��>����)ɖR�����4����X}��}-y�gJ��L0è�,��~��_���4��,�l���]:�Ԝ�?12� M�5��'?���-I5Wv}C�e��b�q��_`�e*ʲ����_��̈́��+U��n��zbAq'E)��R�@��n�9����$��,�e�À)�}a,@e�Y�[;�f?k��� H��ϙ��R�(�v-]�4A��BM�K����͙��tӸ�1�(��y�Kغ�\�B��6�HYQ��'�5l�X�X��<*�
��;,IJS�׸��2*���Z3��3w�
R�N�h�hE�v�De7Pd�K6�I[����O?U<(�$�M�n���}�1Y��$�Ђpscu�Ui_����_i�����s�/?Ԗ$"�1�?G�ӛ3��l6(�k�4��\�2/o^P3���\N>��.u	�~i�m��u��,��_���!�gm�yH0�Mb�k+����<'9�)X�������RR��8L�x�k��o����UtrK�rq�m�����)]�%���r�< �4M:��o.mW���% ��oJ$�JqI@�6���O�y�_g�(H-���{�2_�6
Eٹ�[�����L�-�ڃ��'�iz
�:dM��>8R����꿖��ag��0s���u��z�Ѥ�� "�V:�W�ux�-���&GFx#ϳ��X}s�G<f
��,�+��%Ғ1����� p�X�<*u<=f�]'X�	�DՓ7�gS4�������v�D#8YЩj�]��v=VQ>Z~�a�7G�����8;t�HT����C];L>�S\���W�[�� ��q�ƌ�+�]���L�-&�p�6�����t�D�W�Me��:W�Uu3;��J��QuV>�(v���
�0�5FZ1E���p�ñ��w�"��z�	�2������֛�.��,��3y�$"!lj1�J���	5��s��נs�d��(��i��S��t���-����N\��;�g�ԇ�������<��kr{/����*���ۥhR����U�2���o�$ �X���+� �:T��3Lb(#+��L������]��k��[�J���3��qu�5�k����\h�)�����%����8���e�(�Ȉ�~���uU9��t���C@ÛF���T�L�@�[e��ޏ����@O�N@�-�?UlG�\J �f�R�����?�0���ix˭�J�:f��n�.L�c0M����D����k ����xoZ�	�k&f����g.ڎ����#N}�/��v/d��^��@�ԍ�$��?�};��l����E|ǽ����6d֒��$K}�EI�g���*�q���滜ޞz�,R�e8��(\R���#Xc�E߃ `���6��Go�X8�`j�<F�.=>�0'�<(���R2��W���р��|���X���@�PnQ+<�����&]�`�"I�)�����*���f�=��jE�w#����7]�@�{k���{���i9ʚ@�å��M�	����6�\���8rC���GDBbU�����
APTS[�GdCq�R�"� Y+Й��?�5?<0>�S��kq�BA�l&����LC��X%�;\�ca>���:~�� `#�Ų3��r��08Ǐ�aM��wUd](�P.j��GO(A�f��"��K��}y��\��>�#m4m�Hc�zގo]����/e{£�T����F����n���0r����%��u���A��`�ŗ�Eꉌ~�ɼUc���}�D>������m#4��w���Î�}����0ː0�%����ZwH�����[�BY�C��C�C��~H�T�_�uk�y�=z��(���"���mZ��w�l)���}�>���ΐ��;��=��ˣ�v��,M��YE���%s�*LD�b)?�/Qۃ[�Ǒ�n�p��=�a+u��KK\�4��C�B�yr�лB�!��"e�s��8h����#y6�U�����G�z�JVkDV�H�l��HvrCAv��]ɇ�3��2o�6Ck.3�2.��	�7����B�>�Z����k�����A�=���N�*V���N��&-Y�k�Ó;��BGωHD\�q�&��ȣ�.�&��K�������	���R�{��`�	^Bɇ����L;§V���"A����������z��$���|�/�K� ��{�;���uO,-�=2���ze�Tu1!5�?�4	�G��8�iKA���4K���)��F�:��.�^�#�Y�y���h�z�g���ń���S��֏W���9�>��V󤬂'o3M�ꆑ�#�dH)>��d�IɆ���d־~	i���b?���@�:*��ݾ����^��Jv�Hg�k�����J�mTg���~r)����yȆ��ʙ��-@�Kf_�AZ��E�9`��:�g�c�p�v�P�- ̾���J�~(w�[)t� ��C���1�w!�����R4ż�8��|K��*pPox0��"k��ØS�����V݌Hq� e�_���igv�p��D'��%\�,B��H��&5T)��j뒄r�ՐS��ڿ���5�)��,�#�Y�t|��;"���}�J�fQ�/�_��~є�.��"�
>��d|�Z{M�,)�
V�0tQx�2�������d���`��5��G.��GX0#�XQ5=��r���D��e�Ӽ��T�҆bd�>�����x�9�T�F�㤘��5s�J��FQQ����P$UR̖��T8�ઐ�?��o�岊=�!�I��Tp�e.���Gm׈%Հ��Z�����0Ut�������ÐJ�tМ
��m��,J�`�;}aBJ�)�t���-�CW����P�����Mh��Z��պ;exĩ�D��$M�"X�V����O+[�*�\�ar���AFgxX\x� �ߛ?�6�>����/0�������0p�>��HJL���#���z{�b��������6�M�s�LB}H$Q�YQO�O`�k�^5?┄ ��\���q:��c��L�����xl�Pô��?�(>��ri�MZ��3�<��ӡ*�c0k�a�����Ԉ%����
���}o��S�#��hVzዽ?g�͐o��4ӘG�$H�{Ɖ�]x* 8{1Y������p�A���$���Mu��C?��_�Ǌ�U��-�e|掗�#p"��6��]�L�W�6���AKP�j�s���(T�� ���fT=�|Z��Y��Sg|���*�XW^r���}2bQ`�@�^��X�� E>o�9�T���[�b���Q)y~i��hK1�Y�Oܞ�/d��^̗�BFHU4c3���R���.��liN�-����7{�i<����'yh�#��5��*{-��gv>2�lJ
К��A�{�̯cd
��EN�\R�O��T�} �� ��쿍�Q(n������t�]�$K��͓o0�sG<Y�g���1�:�D���"����������y����q��٣&��X��b���-��Y��� �\�e����������;Y���t-�?T-JA��¡4���c��9�ݻ�T����4ˑ�C�v�6�ٟtv��E�zy�a�e�=��E� 