��/  �
mqm6�w$]�S�VX�:J�#�Zeɒ����7����h!��?VZ�}��rWઇ�]��  ԚS�d�|(Wj)�|Qbr�ۜ�d�
�Ze�5��q*؃|���ye|�|��L}."��2�Hk������t���kJ��Ya�a�
����pg��,�ޟ�p�Q��eгC�Vq�|����D�LDz� _�K2��({�ya�Ko��5�-`FQ��r9������
�r�Ȧa�z�W��T� %��֦ʴ�vb �ǾM���Z3�ĂR�	���ON R��Hq��6�l�誖�,C�LZ,��~�hʙ@Ӯ�p��	ނ��ܪ�p<�u����-����4BEP?�9?[����¯��0�i�,+��(��ByO^��0n^!��X9HxX�)�H�Q='�l$��s7+�,��@-O�*�_��S:l1��~�v��h���
^�Y��� L�7��G�X�G�r��Ê��w O�D�v&4[�/�=�"�@�G��D)7�:_���f�1���zY����/ʌ
�t�4���=�X���������W�y���]M�����5��K�l�ӌ���U}��f�����9�ϼh.x<��V�k�B�� ��d8��fU
�&��PU�0���͊�K�%z "ی7q/eA�w����qj��+��]�E'�6��?�������*��XJ���>�bZX��&@׬'!-~<�H���U��B�8]f���T�ܫ��N�61yL��yn�o'ь"`u���V�7�F+8Rm�U�+2�G�㶳6z�)�R,�tI�r�=�ӓS�ELѨ�����=C,�s�r.�󬡱�q�ފ'3��w�p�?5S6�y�e�T^��F~\$+3j�pO`�� eF|(��k�T`D�0������`�6Z�@�H���lsvk�lMvi&�f}�>� �ϱL����őQ���Q�2��I�q��r�I���8:i7zi�����YSG�kK2�i��_e���?eN8Jꗹ��� l����|���ޏ��8͉#�XtT��ȭj]�e7m�q�����I��<,"� l���]�v��k�Ȑ4��A�'{T���Wc$y���9�?4X���]`NE����ѓ3|��" _������_EiO�%��Ԥ)7� ��d���a��EG2�CG�?T�,@���]���5�\=�pf��ҍ^ޒ�Zn�5W���V�\Hka#]R*7�$�/�K����t�.��nR|�1E�V�	`Ң��Sz�_¿��KV�_k!�����\"TH�e0��Ri`U�Q��
���%=��b��ʴ��E�/���W���+R���&�D�t�^�!�t�B r1@S�DS���gQ��n�V��V�1���j[~[]Z��V��hbn*�Ƹ�3G���$�Lvw��/��������X��963A��m���sϩj��p��9���_�/�,��ġ���
V9v����x[�LI���e��~C3@N&��^W��b�F��6������K*��H�Q��<�r�=�U3
�XV���ﲞS���|�fG!����;�]���Tnڳt��87��_{��-Z��X�u΂�(���w��m��|+�lXԠ�39B4𲱪��LQF�2D�_���bo��H A\N��I����6P��t�D�q)��4�ێV�7����z(]B�%M�~�1<`#��G-A�Zv"�%��X^	+�$4:c�����0܈����|���_�9=L,��Q~���<����]����I��Y�-�<3B��x�rT��BH��1��[�����1�_���Z�{�#<f���`J�:'�w����+������p{��<P�,xb�1`�[	����
qT�(�(O�J2	��]�MM�r�HcIF�|��
��$���N�~Y��G3���(Mc�#b��LqWӻ���f�f*R.�a}�o���x�z#wE m@e�~��ĥ����aTV�C�EF�^J8��6�Uآ����	l�0���&�Q�8�p)�V>�&�T�ݐ`��	���_�������5A<4�)��ĥ[��3��Vw�;E��oS5%|�m(�*�1Kg��	OXnZ;�po?��ںeR3�髗�B�
�R�DO,���<��*���Լ�G%�()n���긟�ht�A��
?O�we#�[�c~N)!ڞ��݆�� �\��^-��r��XZ*VM�2e\�������`pOk�]���u���Xj���$�)��@�3��E�׌��V�=�YY�+cs�\�O�ί-��t�L�N�{N*f@k�H�����!��M�� i�"M��c|e>Iu���r?ɶ�Hw������c�@8�����P$�d!H�ե�3@��}dO��z����%��V;�?��2�B�(s[d���hgZ�¼����z��_uM�dIG^��8iv�d��A�U�5
K�sB�i(m��(�E,�$�D�xԚI�7-��UI��ep����������몫8~�3ϕ~/���~�J�|���9	d-~,��Բ��R�lp����w�^ĒM�ő�V��9��a;��*��Xc����Y~��Mz�X[��J��O����I!��-k� jZ�t&>.B\��e�*��h
��2��.�x��֚�o����+�S�Z�8���CU\�M����偂A�v)�2����{��Q� o�*+v�ʭ�l��.]�.����"�E,A��Nk�3k}%8i�mk�jE��E��N���C�\xz̷}�`v/��*-��&��v˱��L�#�:�8����Ss��x�伬z"?P�%
�0F8�3Z0�n���G\q����bg�1������ΕC��M�&�w��� vU���Rm��f��aV�^�b�J6�9���g�<�� �=��4X�(R�����\� 
��5O�mQ�ma�W#�!�ٝ��GQ��w_�cYw�=�3��w�M��s]����9Kɡ����g_�O�lpQ �m|A<z
3Wy����?%�|���P���K%�2�ų�=��P�"3}>Qc=�d�0�_ �'��a�%D���K�$��ML���s��8��<H�E\$���JqT�N{����xi����]���7�B�+��Ś&먽�qI�M����N�髂d��K��D{=dl��P���ϱ�/݄+~<��KӧΉ�()0'���q�v����5��/��ˋ��{��|Ko[c�v��Y��Z$�D�qh� �ҷ& �O�{]݁2�gպU	�K�ΰ��t�2W �����Ė���3��Q�U�<�ʾ�fJ��SF|�Yc9{eyv��7�_"a�8���������*�D��=;Gv�#Ӧ>��\�+��s�i�d�sA�F�ϗ�+1�oS�EF�>a�	��:����MB�7�11��`�s�'�1��9El��Om��~�T�������B1Tk�5��3,��/�(�L��e����ٺ���x6A�W�m�c�>�ڟM�za���%���NeU3����@��i��S�78:��r�'������%����{�D?DF[���>�YN������b�e��E��������pc��n�aH�]�@n��,�k�e\��n�\FU9h��)a9B&1�i�&Se|���G�Mv���sc�'�:[�&yZ��Ef��p�������oin#-��0�/ �����+��ds�����@4/Kw�,4~�q��I?�=�EEBO��L��k��kv����>x%3�W}�?s��ٜ�����lIF����Y�{3���S�秆���&�H-��Ns�V�q����^d��A�������:����!k��Q���Ir��FAe��|�@���>�`*Ndr)�����5�'@�=u1�	�2E��%o.uKF2�^��n3�3�ac�I��yh�Ӆ�Y�U �B�t�J�ߏ���JifDd�^s�q��r��B��Q����:B��e,^�_k�E��W:POW�����a�|����8o��hz�����3K5�[\�P.�y6�4':�r�Aۇ��un�9��:U[&x��L��D\���>��ӣ#�ь:��U�|!����QIڱ��,�L�q�	�|�W���'~#`��On=��
�y�ܻ�AIj��!/${ݬ]wG�
":2�ւ���:�u��9��S=�Ow���n�Sq�e�ȉq�:�+�"�����,u�k]�ET�"�ȳ��Z��Ŵ���&���V�
8H�ξ¥��Sa"���g��f��u��Y�kt
Eȍ�{q\�(��,��\�\[��N�TOS�n�&�,'y�|�{O�̅4�V�
��� h��!�g]��и[�A.^��`y�����p����>�L�[&���� g^M{���ѣ+����Uc��D�B\a2o�yi��z�#���b!���y�C)�J)g��[1h��2�9c�[F>� �LJ_V�Βߏ�kDTS�=�u�%�����,Eg�ŝ%
�
�JY�&3МP鴾�L����@�LhϱZ�1#�W4�I��r�`)8
y�z���^@�x�'��^�����04l�Y��5$��5�k�ă4&S�9,tUnV����z��T��a�җ�D�*q�t<�Ԗ��`��׾큯֢�v�ET~!����\s�{c�z	n�b�f	OGO�<� �\�|*0�<sk�~[����nY�7���f	[I}m�b�g��@K��Ͱ&h�xB
'۞u 7���>���ï+��bkЊ6N�fwF�}�v�]x��]�տǂA0��{�X����xI�2�p?�,V�e��.��,�D0f�3�}���b�L��QS�n��-4!إj��M>�V (����7���x��ǲyz�������K���i3"
�L)#&m�w]p����J�A�{��۪�v�@(?(�S�҃	 )���"�h! p,�uu0L����0�n�&H����t�]i��NP�y�����a�{�>�}����@q�?�q�GN��E$�j�B�Ш�|�E;a��eʑ��QjId��������L�H����\If墆DvaR?Ƽ�o|p���?�|$$DA�w4O��A,���'�t�|D�+�L2uz9$�k1��h�����R���<Ў4k��xS7Ta�q��u?����&)s\��-aH	|�t>��,66竞yVyn~L�Ӯ�O��tj�\sm�{)�s!X�FH��0��;[��Ԉҿ�!U^5�׌���+�R9W`�X==a����KS�2*���fJ�<.͋s��R��%*D��t�pf��c�3��f�M�sM��U0�kb�k��������oa��ҳ֨v�����2.úfb���pr�6�~��x"Q0QBZ�O�{6Q+�~P�EH�d�U,�v�W�_�=Q�.��{@I��PI����|�a��)��{_Å�"	Y�j��4����g��Fz���|�ۚk����~�p�&�Kά��p�OS�j�yt��MY0ҟ��������薝N���e�S�M�] �*YVbU�{z��m�k&
NW�"�ň�K�1�����'�t_�mD�x��{�hTUl����C������n���%ƞ�?�@������v&Wb��_��cDɁ*c�n�uB�-�
w_	���+�bݕ��4y�"�p,�/��hv'��sƕ����'�+[� ����K���J�c�$g��N�{��+ �H�m�5��Ƙ�)RS�����pjʄ��gS�".4Y�� �GR"�(r��wx�cߪ�z���3� ���<�s�Y���(H��J_֧�rp��v��q�M�%��1����'���q��a܊��b�t!���������P�#�NFK��c������6�7�h�gt���E��������5p�e�zԐƐ��[Tm�3 ������fi�"Y�K`"�Т�H��VEr?���_,0�|�D��xzZ�2�S�	�*�D@[�c��&C�N���USh��V"r taD� g+@��5n����.������ vZ쵄�#�o�I�[�"W	>���g���=��6�2�5G*\��u�`��7���*��	��÷�ߜ�Zg�H;����"K��[N~����l���Ѱuo���7��Hi�Zw�dGC���Spm�e�H���#�B�y��ZslN�'��z���$ڝ�я�����n�2Y����6�[���|���8��4�ujkU�Z��P��a��)}7?�:z:����t\®��{�6�?�v����Q�Xy+�����55i)Q M�i!�Z^@�pt	����oT�sd��9{S���Ax�aP�Ǽ3<1�)�x�l�{�+۔�_��#t*��8�է�p��8��ǞU��+�AX�V�h<�+:���}�ެ\{[*\0,���~��C��<��S(ڌ��ݿ!�u�l(����G�����-�����`UT~[�����臊��oV�zv���~B�OMA����~������vv@dc\ױ�ƻ(��C���j[�3i����c9n0��k^��F����W.�bQ�;ɩUm��$���-�9&[��D7yd�N� J��"��$Y��z�#�#ef����Th["�X�+�=��(���-Zl, ���.?�5_I�����.r@��\[���l����.���1��6�$�3���U�&���:_��m��	�S�o�K�<PR����Ow��Ҡ�W�`<����o ��⦮ᏠځnF#ϸ�z�0s�-7P��yd���@�@B�FV�D��|���Hu��=B�j�h`)���M��9����Қ^{i�OY���^m�0�	�_��?
Q�e��DP7�@#_�-�H6�7� ����{!�8�3-୞�Zi��	[ �m��0a)�S�ק��-줕L�>�o��^���+�To��	-��t�A���bFunah�P¤3�;�욾�+w�tє�1��d�����S)�U�Oe���yg��+\��#���I"��9���Κ[�9W'��Ƀٍ�%��v�	YN��x�^����(MCA6�}9g55U������ˡ�Ʌ��n��Av}�@�6H�N�{�^QQ�'��S������g�{���,5�����᭯7�B?��eWW�4j�s��|&�=�b��b���z�R��MT�ԛ+�X���M�81�q�v.��Q'����2�ٰ?�O��vl��e�[;�T+����oA�_A
&j[:z&�߻��g��qI�/?�$t�����b�j�)b�O{ָd��������n���q{ʦ
��Id���XO�ʇAL��d̉�F��o]3��1|Ϡ�F��f���v��
ֹ��Xœ0[��A��M%}�"(��0�n/ݳU2���u���+�����R4,��)O�����/.�^�!��]����2'^8�Ka��~ �E�|����[;���{��U֏)�JRQ�czR/gU��j��`I(Y&{���-�
�#������jZ?�c��{s9a�ya�}4��aK��ne�Qfd4`��9x�Y�I)?\�~(��EYp�r�@���t��mYzݞ-e��C��Q�p�#1~�i��)�0x��|���_����3S���_��RK)�p7[�������M��*`tH��'R�?�w#�n�����)�Yi�F�WL,��0�K<�jh�1�ȅ��߈݀I������"���q������?��3����V�m�d}v9��hOD�!�59
�ߓ!R�d w>��͗э������X����e/]�ز]��/�v^���������X��{�S�>���OJ	�s���m4�l�p_q�*���c�e���L�9]���F����lx8��ĺ�[�*�1���
�{ �o�{����/�[L�훁r~N�s����8��Am�
�`��A}�`�.����c |# 
=.����C��I�7��q�>Ca�N��z���br\+��T�z#=y8�G˭�L��	�\"��ğ�6��`^s�W�	�!�"X��h�7�k����$�y7���<,���|w����� +�C'��D��kۮX�[��}��m���Χ�c<L�o'�����>�b�i�������o�N��^��a��?���~팷>��X"@,�0���,��@0	�#�w.�_��r}ÞS��)NV+� �7&M���k�H�/��H	%�ǌA0�x0�Ӑr>���\g���;���׳p<|��mt���C,S,پ-v��h��r$9.zT��Y�(H�2��6b�bW@ T����qlK$�.�wg��J�Z�׈ �u���eUJ*Y]�͔��s�w��x2
́P�q�������I�ǒ"��
#v�sTN�4> ���qcY3�?�t���G��)��8�����:�m�F�2��ڝ�F�,|-z���/#F��:y_���&ZQ��C@''_.%D6Q:��kg��B#H���}E����"2Y�E�����"��v��D��R�/K�"z�|*9	'��և�����J*t��y8.,!_�C��h%���{H2-!ZI�& ��p�:�.0��l�A{�yCn�����Q�U��5�Jr����UT�E�:�/�U�N���]"�rj�֦�`��HZǻ���~S]tG,�߸u�0l[�lc�ղ�K�k��M�8���vN�n�2C(�u�����K�~����� ~Z��Kò������������@�I ��UF���̾��,h�`5�C4���f���״ó��YGS|]��)�9(@+�/�x�'c�`����߁���Joryp��P�i��8:�_s �w���~��Pq�ܤ7��Mn���DRi� �<�m2|q��v�I2�^Ƕ +i��P�?�l�,H*���U)����<E�C��u�����ʽ
h8�.84B��-�����'[�ʡ�ʼ4��]G	�u~��c�t�:�j���Д���"��T���%�/�f�m�Q����z�;q����:�ds��P���\J����⣰�!�����\�x�����|w&�ҵ(����ԝ�n�ṗLkf8��;Mq�A�vF�����()�� 9�}�`�=B����"ˈ_y�8���?��6�^���@���Z_-���:��������R�#�