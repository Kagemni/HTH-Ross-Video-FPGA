��/  �^���H�Ҭл΋2;�9�i���t9"j�i�z3]G��`����$[X:��5gn��o=��Q��E��l�w�p�/��ag�I<����V��33<=r7V&��1?�~�M�#���b*=��Db_?���v>���D�!E:	z!�IZlW�0jA,�M��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n��:>7ߎ��Ғa��H�Ɯyї^sXz�1>l��^OɧF�e\p��.�Բ�O�mVZY�5F��6��Ѕ@?�;.�8Il��{�mp2�"f=���Y K,�J�T!a�g�Xp����6q@A\2�J��,�JR�	�d"��������ॳW?E��I�����wF��q����7'��ve��f�+��(��O��C|t�or��vP�	"t���kk�= >�,�C�%DG�  �j��K�s3d�at��<�d#�g��8ӥe��~�Aqg���1EJ�yF�\�����˄���1��ՂƎ�_z�1y��ζa���CW<~H�-4�9x/�e���~���S?gl����b�76j�� ���'��y|�S�N���z|7�U���nlM�H�UT���gp|�w��B7�K�C��|�>��G"��������X`P��T�m��ksC���t�794�w{�qhN��̬%��K���0w��.�bT������� HTEǟ(6?8�[�S���; <}��c�W��'U�ؒ���aH����f���������V���mK�j�u�������J^�ҝ�{�OK��-��Ug��f%�ŝ��c�Sy�"ٞ��˥�&\C��ψ��b�>�5����[����O-��l23��y)��>�8ŭ���9��$�i9��x`X�F]Ǝ����i�7�pr�� �ZWw��p�� .՟ꤓKɢ���GsI�����3�O��Ta���r�=(�ƃΒ�׶y��A!�ǚR�}���Ϊm�G�� ����=l�o���LZ���
D��X�}���2"�.ˉ�N���Й���LP/7d+C�Р#~�RɌ�8���ą�m 
�k���H8U�xa�4�Ya��03�n�܇T9�
��!��޽W!O�NLy_�~�v��kY�!������6�iă+!�ס�i�<6�yV�J�*�	�\�H�W�|�x̭�.ƾ����[���s+�G�9�ΰ%q��R�'���"��șpT���RL����;�J�c��pX�m��# %�Fg@���Ú9�����ӫޗ�.j3��6/�N��p���B41��|�4����q�eQ��'��}����U�wd7�,5h�����:G�MC����!?��)�XXZ$mmBx�=G�
�jPb�ߩJ.�U�C%x�IVg4d�Z�!���4���7��G?����&�V�N^���N�먽�zB�0fo���k����F�H:����pA���y|;ʗ(����Tݓ�[����"�~7��t#g���g��(�Q�@����=|P�	�����T3���T�1�g*�YJi�����W�Q5|�|nJ��*C�\'�!�	!uӜ�&����=�mu���!�
�Y�S�����əb�� o#O��������%�| 2g�;&��՟�R���ř!�/o �N;�Q]`�N��1�j,��������ľ#�]�
_9ؑ_4+ӿ�;%�Oqj�C�`�N�k�?������jD���`6��)�V��Y�'��`<�g�V�����(A�UO����_T��0�*��3�{�4�����]ر��"�]Ia��J>�i�Ⱦ�*p�K�6�2VSHy���N>��ə�m�8<�j��w>���ܝ9{?��o�7�J���}������(¢��Lp4 k�H0"����-�aT�m��z]�|�y�]H
<��h��ƶ�s�"2�5�>�7V��D3�<ҷs Q^�6�T��=i����{�h�uO>���WH�ػ�XwRgR�\�lz�H��K���3��9j�w�ţJ|�+�2��!�ԇ�x)���+��3�z�U�t�s�p�R��X�E�/��8�f�%�G�>��R6a��WrM=��T�Y����(����#q��4�F�F�|eY����8Z8�Z�MM��'�#�Q��%e2��쫟��e "�E�r�#����*^<�&���D�������Z�g��q����J��Ѩ���r�b>15��4hz-o�f����#�"��\�)��-�]"N�:�&
UP��0��+#g�<���K�d!-�CP���L8�����5<ac~7�4�9xT��QssΧ���&�wbk cw�����X��KH�%2ʥ*p
݃.2I����>V#=�q�z]��ׅ�z����6=�@�>ŰJȦq����)<��s�)q�YJ�gQ�LJ��9��4���a�>ٖ�|�E���!�lEv��\��yip�Gd�F�ԏ���?���	�<ޫ*3�n.�KZ(��ha�$�*����.'@��36�z�LS��<����2De��q��78�]�=�=�@l�;c�Vб\`�{�
iL�r��I#0�`n>UcLGm��0�������q�:��z��`C�k'��>$�ID�������iA�ׁ�3�������Ŵ���	��}�5��J�]���%�-t$��Ս��i��]S��N��7�Ho	���ҳ7���ȅ��	��.��:>���=���gk�Y<e�z����@�O�)�A���{�3�.1��74j��B0�@��Is����~��*B�x},rU�%{�diH��Ԕ���Q�Q�|0���3�.\! G��y!\	75K�X,����/�Q,H��h���mn�9G�آ��[8ԇwL�������wv�Rj�ܗl��.>�-FOCV�8S��Q�3�P:���
��z��_Ї?YK��.\��B�<e�f��@�n�3ܣ�u�N�Ơ�+ƙ0�:pC��
������?r6��/�_��B��F͇]�R�9'oBZv�X��6?n����Kp�����	ׅ,��Ru�y���;N�%�H��u�7��S<y*|*�)��I�e��-@��:Z�Y+��Uy�'��|d�����N\�7����	����`�Ia�Ue?��`��q3O2��ᰴ�7�i'I���'��~���lşJ`�7%v�z�ϖ��t�p�S�T��v����w������И�/�p%�"H�jg�SXt�J�Q�_��!������w�T��Q��'���b,&Y^0cW���:?k��=�ӦO ̲4ߥ4���
��4;f�;a5[�{2��B���'o� ute֕+5���P��P ݢ�����]VQ��[`�A�6OR,Hc���n��,u<�n�F6��0�e�؞���@��u�r�S�����I���/�pbC��wE���"n���]\���k�̰����s�`ۓ%�h@��N�G�r��_9'��^��!�Ī5d!�Qp������e_��)��V�}ɐi4��d�$�&�XE�A�q�^H�B����u��R��wi}?�ə���%R�^׉2*�:ǁ��-��	h)F�ٯ�@�f���\Ο��L3=��)Q�(��=iB�l� ��c��ix$��h71b�E�q�����R��|w�hj�m�;����S]�/���yn|��)AJ�]�t�����x���d���������,�6��u�tψ�Zok�o�@��أ�v�u0��6� ��=L��F�0|�w7]�9s����q@l�m>�l�*?��x���H~�?f��\hP�~ k�!��x���9$�ϐ:���T�5�o���w���EXVM���	�ՊSa@���;�vD��u�T��@y[�[ȚPx�����:$"}T��U�{��_�Z^��B�?�Z��.L��d����b�]L��ӣN$�r'��ʪ\K(�n�e�k�Q*N�Z�j�H\!)L��`I����Lr���
�ҥ�1�����:w�s���CeB��I#�>v��JS��f�#� ����/]�#IT��\�I�ѱU
��$�;N�c���]�T���`7���s��<{����[�advHq@�A9��g9�M�r��Ҳ��X;��/��=ފ�cY�$���L�5��V��`���!7S��>���!���H�9�_;�������r�|��㉌�^tR�M�~��Jm���|���pT�sǝ�8!��["cs�)N
�J#�I����ָ#ҧ�M(����@߱x$V���Y�$��D=�0ح%��/�����,�r��������n��U��$x}�{�{��p�7;���H��񼭢�բM�Z����(q�-� ����,�n��~�y�w9�i����=F�����&r=��R`Y�ڭ[G����޾���YUNAQ��dʆ@|���2DM~J�
LCX'������3�B��|U>�7�Dp�����F-�g�Ŭ�̲�}�+��D�v�լ.4�l�s;<�r���z��{t��m&�'�ͬQƃgDӊ�WY�!��F~�AJT���}���h<i�����Hk^ؔ�����	�"�����Wx�t/ҙ��I0��1�?�|��[�ZZ���+h�����Z���^Z�<Ha����5�!��F���B��x�����2�Y���5��8��)z�	\oR4�mi��h�z�&�����XpX	�-+���C�U�,�*�'���AD�8%�̭�+ M���>N�`'_2�zL6��sU����H�Y�O8�o��O���ōf=��ZuA�������=SQ����we�Ï�bu<��}c����W�(��Pn^w�IuB����"b��:��?��~ݫ�b�g���bp�����P1����1
s���>7(��'d�t	%a�h��bS�R����_Ng���Ƥ=A��j�{1э�>��D{iR������^y'v��чN�$�A���j���A�� ��]���0 dB�>��^~��߉�H���_����>:7,���9�h��3����l+�+b�j��ӱs��Qf,���.I�ˉ����sT�pX�}˃��R�OF�׷��<����M��zK8_z\
f[�3j����I^��^M/�3�%YB�7� �~�W��V�jK�f��DV:h⒋˵�X�k�O3��m����;��I���L��Q=C����{��*���x�Z{$qf�Ќ�A?�D^��,ט�K�6MԵR���]��ͲR���9�a���+��<���6��s���j  �)�����:A���zU�og���cZ\�3f�06�14z,�/C{5�n-:;�-Rz�}�\4��<N�vjHFQ�92��y�	$���H���^�q'���__L���q/w?�j�R�NP���jg��}��Ƿ�=�]�I�d�pX�L� �~J�
��u����q���`|��9��Lt��Nw2���X����k�f9����y�>�P���M�����GpxI����7`��Z�<������ע����t�����������Aڲ�=�ڛ��Ȳ��&H���*Y�n���Zw!n���y���]v��A���4��(	�tf��9�VE�M?A�xL�?�i��������s���r�xF�	4}$D��q��(C��pe\o=b�-��������fZ�ٰ��E7�Iv��ⱶ$֛�Z$�Ko����(R$A�G���aN($��`��x�w�"�؎H��v�Ĩ]0o�7S��=� L*�!��ͧ����� Ҵ�W���胁$���|O 1