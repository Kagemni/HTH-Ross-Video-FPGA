��/  �/�V��6ܼ�� �'J\#v���>B��G��%_�!���G��6���߲ìj6�GE�kPN:�{��!u"����vw�����k�p�,�f�V-�#�sV�[��T��\���4�+��G��os�|>o�D]L��x�9>���TQ-��h2ũ��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n����D3ӡ���p"�pM�x �GIc�W�	� ��S�w��Jƙ�����O�A|$a?<2�9����g���d#X[~&/Y�J�> -4���}Kȟ�U@��[�)�S���W�Oq��>�n;�/�§Ô-e���RS�/��`z�����F�����D>��O���c}��i�L~������q��Y�M�&�����g-f��B˼#\/%�)��U����g8�¨,�x�5T�#@�VH��OM"� ��a�ab��:��~��	[!L�r�~��^�'�����6���R��]�X"�YFJ�I��@Efp�[Ԣؒ���N�na�b�����	���q��׈���#�RJHm�|�I/cܾ��.
ޖ�Q��j����Y-̋���@��=\�K?c����C�-!om3A!�pX���'A	zT���-�� 4�Q0�D	!���b*;��C~�V���s��,q�<`�JJ6"����W�w���)��cg�dҐ���D�JR�n�'Cg��#ml:&�����C�MP���m'���D*��a�'~�៌�B�P�U�%ih�ӘV >�do�BS�'@�'�����	� �_�+����(�;�QOT�X�P#�%��ћ�u�U595���,��0��I%d��лIc�V�u1��<f?���F��s�8���L�:$����j�ھ�Ӱ0p{^��t@��"X*�&���t�%�4��b;�Oȴ�as׉s��ۋ�N��}����]��}ށ�����2�Nn����K�}ǣd�xz�z����fbgT2�n:��s���8��_�ŧ!Ղ��s��)�Q�%홓�ΪA-�Ƴ��~�X�{�������}S�U�����T�z�nk�>:aV�[X�����֊�" 劍�ʝU�\.�R����U�q�9�ѥ�0��| �RN�8k�,��q�#	�M	�X3(��!�	qr��$�!�5��D��QS�� ����W�#ndDF�ަg��<�$�R�+�a�j�{N�鈩��$�d�PGv��f�-!�0ST�y,����H��7�؞�3�<Z|z��o0�9ʐ�4�߬��;��V1r\6��R�T��Lq4�b�6��Hn��0�1L�to���}�4�2��{jᇨʁPǪ�,s���\���}4�����p.9~2����sgK�Ŧ�T��?��4W�6QHܫ6�d����Y��=�:�o"�<c�0jo�為9M�O�[��*[�չ7kz����ޥ`����̈́J+�I!��ke��h�m:O�lʕ�j�3,���+ճS���ùg�t(��"��Ņ�����(� ��+#��'xN{�Lj?^�X
]�W�-	9��F�r*޾l�mԻ{n�O���;ii��Ɔ����SMP����D2�v"4%_�6��\ޚ=NV�!lT~&���y*��?4�i;�*�[�6R�>M��e$�m�����������BjM�ĎoMD|"U��*.1N�#�O �K�����B�O/��m��f��lM��ȲU�hV��[����L �?�$�RV�s Y~���eXD*r�E~q~�N|1���Ȳ�Џx䗲;��W���bq{c�{$�`��Y|�V\��jm[��o,�r�9]AJ%JZ*����6>�w��Z�PW��V���v/�f�}k\öU�<�\��:u��yR�1��VҮ�IsZv:�?J���d����y��#Gy�G�6,�~E��R�■T���j�'a�'�7� ���U|[�ܽ���L�C�y�����~N�Ei���ɖ��!1'�u�`L1��#7Q0�M�	��Djy��*W)�. �on�y��9���m6h� y�Fƴ
�+�kL�=�[E&�!����=l���֣��"^?BaK6JA���������n�e`�Ty5q�+�\ܐ��h�YX㔀�ѐz������?}���?�k/g�Ƞ��V�@IZ�!)+�W����$��э�Q�����Dω�cE꒻�b��Z���b�'��[�d���ཾɅd�����xv�穙�d���:V���e(��6s�
�mQ�:�y}S���iM��0����r�����n��KV!"ߌ�fg�q��/c:e����ʨ�OwZ���7u�,��\�A{�B&�w���ȬL �T��N�1�1?|ߋJDD����su������⋈�!�U|�j�^���,hI���=d:��!���u5��|.����!���Lc1;�Y��Q�n��Э��
�s'��v���3�f��0c�;���t%1��O�#�+':��4#�����cR�\`5�0.$�`���l��F���\e��a
B=�1�y7.�-��à�%'`�� %\Ջ�=��=�a�ܭ+V|�g�������`��%�kF��,� \W����]���