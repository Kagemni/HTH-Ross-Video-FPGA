��/  yR��Sc��V���L�8���.Aϡ��g�]��)t�rJ�3t"���	�<�<���༟�x�9��t���Yx�j*���7TN�|�a٦wZk|Z*2u��!)��9t_�L�YU*!_m�K� `�e��p��B�[A̓�4aMZl�_D;N�nQ�d^L};��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n�W��ߌN��5=�8�:N|���gp�P�ظ��U��)�& g�J����[��kC���Rm0�@>��$9P$[��k�jm�Fv
�>v9Z��{�#%"0�k��<p7�#?@�mO/ �w�t���w�⾒�Y��A�����k��^DX�D�3?���{S�+9��0�M�(�98�oL,�zwR점�tp��� J:8k�/ĥ�U]�bO��V?=��:�mڜ>UAgk�j
�����:_�k�MҩQn��g:r_��=S����\��do���[���U�z�� B5Ť��Em����R���.�j��c���q��Ç��Q�.��ڐ�fi��L�2V�CC���Fƀ��(s:��Q��V�3ְ��
H�d; �!Ł�*��u���V�����B��wp{PA��.暒*�0����g�jpb>~y����w+����ӡ���kA�}#�]���iY��͐�:���-b�0`Q�k
|'�G�&70�MXƣ.�7�/F�-��e@��l#���v���Kw��q�,E�6o�{���?�
��J�=s����t6$�l���7��E�?��"H���)b&3a�fa�?�6���ܮ��j�ٟL�yf5A7�&����xG�����"�ث`���'n�Ǯ�"W���Q�ʉ��8���֥�~��=�J蛊`I�Y���N�p�EAo��\�Bva���Z^b��6��I�=��'�N~�>O)%�ͱ����Tfi���W��4,X�,�S�S������0��%b!��ۜ#�'��ށ2���:jA$.�uFdS�� W���j=�B�c��1Z��B�s�����n驘V��X�L�ls�*C&k �TZ����v��W6»�1����YV"pg_�b����}��Y^�Ex�tφ).�>�k���
�a�B�U!�nG�}�na�[�(	�}�-�P��(M���vR"��1K����KuN�0-9{!�/��=���u7��b�q1R��(k�Hr'> �;eB�o�sR�n������=m��ő���d��s��DVu�F:"�&S-���br��o$��9�����>][̪�K��n��R��lc�Qe�1�����l��<�Xg�U�Ӂ~�*-�4�#t�hl���Z��=/�r|"��%jt{�(%+�=��k��4������}�Y�8���O����V��,0r��z�����J���� ?a]*|�%cY7v�����d�oU���|������keD�E .��&̜���FD����jJ�1��� b ��U�5P9j"</G	�r�7�[����� b&i+���>g^gI;��v�ٜ>�D#�76�24:8����ĝ�4s�m];����;v!�H#�_H_�Cg�4�RKy�X~򹔬^6g�<x?�}���V%y���K�[��-EmTJ��<�$�Z�v>��I�����}kt�Wj��2��?-�qҳ�fD