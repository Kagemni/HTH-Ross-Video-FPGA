��/  ��:�x�]<�`��!R6k�S7	(�)���7`.�kA�}���}���l��^���=��3F#��M敢���К�[J�E���r���R��6"��KU|ȹ�'�_�L"�xC}_�;8T!3C߻(pЌ��G�����}6��\��i�=�7��7z��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n����D3ӡ���p"�pM�x �GIc�W�	� ��S�w��Jƙ�����O�A|$aC����e4P!c�O��|%)��ve�.>qG��QܳG{ρ�V�+z8�;[��KM�[	�$G��x/�����8W��m��9�@[�&�!8s�� j�vsJ���è�R�p��@L���(n��&)���8��m%2:��"Ga+�}��E^���٣�0�Dύt@���e�b$�A��U��F�D�cڮ6�����w�W"�|V@U_��V��Ά����78�l�Hd�j̒7���w,��������p�x�[���B�=�:�^UF٩�h�ײ
J���Q�����"F�W�pΝ(%�K^`B��uS��2d^>���z�@�~(�m�"��?/�,���b�L��V�>W���G����M����yG� �,"���[��c�o�ʈ��J=o(���>�+�i�zMނ
2�nfu��n&Qͪ��;?�!?�gb�f��d}��2�-��6���6dwP%d��*�D���=w��c��qUj��k)5˃�����j|W���}���]�s�]$S��0������@�n�kp��\�."���u�{��j�B�X�PCk�I}�%��v�B/)_���/Ԍ�_T��@��ٺ��<�|�+��5dH�	\UM;�W�Iw
�P:Q|�m��)����2kرU��;��g�o��b(��"Mi����ݿ@m��Dϝ$p�����|Z�0�����3�H*��K���Xt��$��%�����D�G9b9������uB��j�j�8A�}�o&k(^��c�oE�T�y|˵�u�=��\xJ9�ɗz
�e�ٯ���{aD|�B�9
�cd#��w�-~��|��pm��}�,�KgN-�ѨP]����y��<�[���x��T׆,Q�id��R�����Y�.�{��Q�C��x��;],lXS��|F,�����	:�gU�qβaf)%�;�ʂ:1tFٲD�ru�Gز�%�6�n���˧(�W�,�#-Aqdf[ܯ���|K�;����>h�����|h�laOwO&�9X�ӰԌ�ck����[a�"���K�'�2�w��dR'�m��E�fIu$�e� ���M���66��I�t��.���J	�����yl����M�E�&��)�EC����ŋ�''/EM'�$��鹩�<s8�L�PLgN`����Ɗk�1�QKX5�J�}�*����cM_�:��v)����1��E�z,{5Cګ���(�T�Q��>;T7���6�ڨ�߄��S�u�k5�������3kQ�]��K$)@
��B�'Y��/1a��)�w%A��2�����p,Ǵ�-��f��eD�!&c�{�@�d��wm?�#���[>��/����r��yT�?WÛc�h�}CF����{���s.d�[D�>�w�S-(4όZ	�y%�bL�Ƹ���i�e)lC�d��1]@��w�\��A(�mf'lv��V��"q��Xu8�E|;�klJs�)��i�Z��x �+{�0�@}U��Ga`h��;<���v��$���|"u#�1M:�66(�i���4���F�����C!s�cͷ4;�K�S�IB�����R�c�<|:�ߧ#v�䝽�#2h��� ���j^a����ux��=Eu�%��消���k�'�