// s5_iob_sdi_tx.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module s5_iob_sdi_tx (
		input  wire [0:0]   pll_powerdown_pll_powerdown,           //      pll_powerdown.pll_powerdown
		input  wire [0:0]   pll_select_pll_select,                 //         pll_select.pll_select
		output wire [91:0]  reconfig_from_xcvr_reconfig_from_xcvr, // reconfig_from_xcvr.reconfig_from_xcvr
		input  wire [139:0] reconfig_to_xcvr_reconfig_to_xcvr,     //   reconfig_to_xcvr.reconfig_to_xcvr
		output wire [0:0]   tx_10g_clkout_tx_10g_clkout,           //      tx_10g_clkout.tx_10g_clkout
		input  wire [8:0]   tx_10g_control_tx_10g_control,         //     tx_10g_control.tx_10g_control
		input  wire [0:0]   tx_10g_coreclkin_tx_10g_coreclkin,     //   tx_10g_coreclkin.tx_10g_coreclkin
		input  wire [0:0]   tx_10g_data_valid_tx_10g_data_valid,   //  tx_10g_data_valid.tx_10g_data_valid
		input  wire         tx_clock_clk,                          //           tx_clock.clk
		input  wire [63:0]  tx_parallel_data_tx_parallel_data,     //   tx_parallel_data.tx_parallel_data
		input  wire [0:0]   tx_pll_refclk_tx_pll_refclk,           //      tx_pll_refclk.tx_pll_refclk
		output wire [0:0]   tx_ready_tx_ready,                     //           tx_ready.tx_ready
		input  wire         tx_reset_reset,                        //           tx_reset.reset
		output wire [0:0]   tx_serial_data_tx_serial_data          //     tx_serial_data.tx_serial_data
	);

	wire  [0:0] xcvr_native_avgz_0_pll_locked_pll_locked;              // xcvr_native_avgz_0:pll_locked -> xcvr_reset_control_tx:pll_locked
	wire  [0:0] xcvr_reset_control_tx_tx_analogreset_tx_analogreset;   // xcvr_reset_control_tx:tx_analogreset -> xcvr_native_avgz_0:tx_analogreset
	wire  [0:0] xcvr_native_avgz_0_tx_cal_busy_tx_cal_busy;            // xcvr_native_avgz_0:tx_cal_busy -> xcvr_reset_control_tx:tx_cal_busy
	wire  [0:0] xcvr_reset_control_tx_tx_digitalreset_tx_digitalreset; // xcvr_reset_control_tx:tx_digitalreset -> xcvr_native_avgz_0:tx_digitalreset

	altera_xcvr_native_sv #(
		.tx_enable                       (1),
		.rx_enable                       (0),
		.enable_std                      (0),
		.enable_teng                     (1),
		.data_path_select                ("10G"),
		.channels                        (1),
		.bonded_mode                     ("non_bonded"),
		.data_rate                       ("11880 Mbps"),
		.pma_width                       (40),
		.tx_pma_clk_div                  (1),
		.tx_pma_txdetectrx_ctrl          (0),
		.pll_reconfig_enable             (0),
		.pll_external_enable             (0),
		.pll_data_rate                   ("11880 Mbps"),
		.pll_type                        ("ATX"),
		.pll_network_select              ("x1"),
		.plls                            (1),
		.pll_select                      (0),
		.pll_refclk_cnt                  (1),
		.pll_refclk_select               ("0"),
		.pll_refclk_freq                 ("148.5 MHz"),
		.pll_feedback_path               ("internal"),
		.cdr_reconfig_enable             (0),
		.cdr_refclk_cnt                  (1),
		.cdr_refclk_select               (0),
		.cdr_refclk_freq                 ("148.5 MHz"),
		.rx_ppm_detect_threshold         ("1000"),
		.rx_clkslip_enable               (1),
		.std_protocol_hint               ("basic"),
		.std_pcs_pma_width               (10),
		.std_low_latency_bypass_enable   (0),
		.std_tx_pcfifo_mode              ("low_latency"),
		.std_rx_pcfifo_mode              ("low_latency"),
		.std_rx_byte_order_enable        (0),
		.std_rx_byte_order_mode          ("manual"),
		.std_rx_byte_order_width         (10),
		.std_rx_byte_order_symbol_count  (1),
		.std_rx_byte_order_pattern       ("0"),
		.std_rx_byte_order_pad           ("0"),
		.std_tx_byte_ser_enable          (0),
		.std_rx_byte_deser_enable        (0),
		.std_tx_8b10b_enable             (0),
		.std_tx_8b10b_disp_ctrl_enable   (0),
		.std_rx_8b10b_enable             (0),
		.std_rx_rmfifo_enable            (0),
		.std_rx_rmfifo_pattern_p         ("00000"),
		.std_rx_rmfifo_pattern_n         ("00000"),
		.std_tx_bitslip_enable           (0),
		.std_rx_word_aligner_mode        ("bit_slip"),
		.std_rx_word_aligner_pattern_len (7),
		.std_rx_word_aligner_pattern     ("0000000000"),
		.std_rx_word_aligner_rknumber    (3),
		.std_rx_word_aligner_renumber    (3),
		.std_rx_word_aligner_rgnumber    (3),
		.std_rx_run_length_val           (31),
		.std_tx_bitrev_enable            (0),
		.std_rx_bitrev_enable            (0),
		.std_tx_byterev_enable           (0),
		.std_rx_byterev_enable           (0),
		.std_tx_polinv_enable            (0),
		.std_rx_polinv_enable            (0),
		.teng_protocol_hint              ("basic"),
		.teng_pcs_pma_width              (40),
		.teng_pld_pcs_width              (40),
		.teng_txfifo_mode                ("phase_comp"),
		.teng_txfifo_full                (31),
		.teng_txfifo_empty               (0),
		.teng_txfifo_pfull               (23),
		.teng_txfifo_pempty              (2),
		.teng_rxfifo_mode                ("phase_comp"),
		.teng_rxfifo_full                (31),
		.teng_rxfifo_empty               (0),
		.teng_rxfifo_pfull               (23),
		.teng_rxfifo_pempty              (2),
		.teng_rxfifo_align_del           (0),
		.teng_rxfifo_control_del         (0),
		.teng_tx_frmgen_enable           (0),
		.teng_tx_frmgen_user_length      (2048),
		.teng_tx_frmgen_burst_enable     (0),
		.teng_rx_frmsync_enable          (0),
		.teng_rx_frmsync_user_length     (2048),
		.teng_frmgensync_diag_word       ("6400000000000000"),
		.teng_frmgensync_scrm_word       ("2800000000000000"),
		.teng_frmgensync_skip_word       ("1e1e1e1e1e1e1e1e"),
		.teng_frmgensync_sync_word       ("78f678f678f678f6"),
		.teng_tx_sh_err                  (0),
		.teng_tx_crcgen_enable           (0),
		.teng_rx_crcchk_enable           (0),
		.teng_tx_64b66b_enable           (0),
		.teng_rx_64b66b_enable           (0),
		.teng_tx_scram_enable            (0),
		.teng_tx_scram_user_seed         ("000000000000000"),
		.teng_rx_descram_enable          (0),
		.teng_tx_dispgen_enable          (0),
		.teng_rx_dispchk_enable          (0),
		.teng_rx_blksync_enable          (0),
		.teng_tx_polinv_enable           (0),
		.teng_tx_bitslip_enable          (0),
		.teng_rx_polinv_enable           (0),
		.teng_rx_bitslip_enable          (0)
	) xcvr_native_avgz_0 (
		.pll_powerdown             (pll_powerdown_pll_powerdown),                                                          //      pll_powerdown.pll_powerdown
		.tx_analogreset            (xcvr_reset_control_tx_tx_analogreset_tx_analogreset),                                  //     tx_analogreset.tx_analogreset
		.tx_digitalreset           (xcvr_reset_control_tx_tx_digitalreset_tx_digitalreset),                                //    tx_digitalreset.tx_digitalreset
		.tx_pll_refclk             (tx_pll_refclk_tx_pll_refclk),                                                          //      tx_pll_refclk.tx_pll_refclk
		.tx_serial_data            (tx_serial_data_tx_serial_data),                                                        //     tx_serial_data.tx_serial_data
		.pll_locked                (xcvr_native_avgz_0_pll_locked_pll_locked),                                             //         pll_locked.pll_locked
		.tx_parallel_data          (tx_parallel_data_tx_parallel_data),                                                    //   tx_parallel_data.tx_parallel_data
		.tx_10g_coreclkin          (tx_10g_coreclkin_tx_10g_coreclkin),                                                    //   tx_10g_coreclkin.tx_10g_coreclkin
		.tx_10g_clkout             (tx_10g_clkout_tx_10g_clkout),                                                          //      tx_10g_clkout.tx_10g_clkout
		.tx_10g_control            (tx_10g_control_tx_10g_control),                                                        //     tx_10g_control.tx_10g_control
		.tx_10g_data_valid         (tx_10g_data_valid_tx_10g_data_valid),                                                  //  tx_10g_data_valid.tx_10g_data_valid
		.tx_cal_busy               (xcvr_native_avgz_0_tx_cal_busy_tx_cal_busy),                                           //        tx_cal_busy.tx_cal_busy
		.reconfig_to_xcvr          (reconfig_to_xcvr_reconfig_to_xcvr),                                                    //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (reconfig_from_xcvr_reconfig_from_xcvr),                                                // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_pma_clkout             (),                                                                                     //        (terminated)
		.tx_pma_pclk               (),                                                                                     //        (terminated)
		.tx_pma_parallel_data      (80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.ext_pll_clk               (1'b0),                                                                                 //        (terminated)
		.rx_analogreset            (1'b0),                                                                                 //        (terminated)
		.rx_digitalreset           (1'b0),                                                                                 //        (terminated)
		.rx_cdr_refclk             (1'b0),                                                                                 //        (terminated)
		.rx_pma_clkout             (),                                                                                     //        (terminated)
		.rx_pma_pclk               (),                                                                                     //        (terminated)
		.rx_serial_data            (1'b0),                                                                                 //        (terminated)
		.rx_pma_parallel_data      (),                                                                                     //        (terminated)
		.rx_clkslip                (1'b0),                                                                                 //        (terminated)
		.rx_clklow                 (),                                                                                     //        (terminated)
		.rx_fref                   (),                                                                                     //        (terminated)
		.rx_set_locktodata         (1'b0),                                                                                 //        (terminated)
		.rx_set_locktoref          (1'b0),                                                                                 //        (terminated)
		.rx_is_lockedtoref         (),                                                                                     //        (terminated)
		.rx_is_lockedtodata        (),                                                                                     //        (terminated)
		.rx_seriallpbken           (1'b0),                                                                                 //        (terminated)
		.rx_signaldetect           (),                                                                                     //        (terminated)
		.rx_pma_qpipulldn          (1'b0),                                                                                 //        (terminated)
		.tx_pma_qpipullup          (1'b0),                                                                                 //        (terminated)
		.tx_pma_qpipulldn          (1'b0),                                                                                 //        (terminated)
		.tx_pma_txdetectrx         (1'b0),                                                                                 //        (terminated)
		.tx_pma_rxfound            (),                                                                                     //        (terminated)
		.rx_parallel_data          (),                                                                                     //        (terminated)
		.tx_std_coreclkin          (1'b0),                                                                                 //        (terminated)
		.rx_std_coreclkin          (1'b0),                                                                                 //        (terminated)
		.tx_std_clkout             (),                                                                                     //        (terminated)
		.rx_std_clkout             (),                                                                                     //        (terminated)
		.rx_std_prbs_done          (),                                                                                     //        (terminated)
		.rx_std_prbs_err           (),                                                                                     //        (terminated)
		.tx_std_pcfifo_full        (),                                                                                     //        (terminated)
		.tx_std_pcfifo_empty       (),                                                                                     //        (terminated)
		.rx_std_pcfifo_full        (),                                                                                     //        (terminated)
		.rx_std_pcfifo_empty       (),                                                                                     //        (terminated)
		.rx_std_byteorder_ena      (1'b0),                                                                                 //        (terminated)
		.rx_std_byteorder_flag     (),                                                                                     //        (terminated)
		.rx_std_rmfifo_full        (),                                                                                     //        (terminated)
		.rx_std_rmfifo_empty       (),                                                                                     //        (terminated)
		.rx_std_wa_patternalign    (1'b0),                                                                                 //        (terminated)
		.rx_std_wa_a1a2size        (1'b0),                                                                                 //        (terminated)
		.tx_std_bitslipboundarysel (5'b00000),                                                                             //        (terminated)
		.rx_std_bitslipboundarysel (),                                                                                     //        (terminated)
		.rx_std_bitslip            (1'b0),                                                                                 //        (terminated)
		.rx_std_runlength_err      (),                                                                                     //        (terminated)
		.rx_std_bitrev_ena         (1'b0),                                                                                 //        (terminated)
		.rx_std_byterev_ena        (1'b0),                                                                                 //        (terminated)
		.tx_std_polinv             (1'b0),                                                                                 //        (terminated)
		.rx_std_polinv             (1'b0),                                                                                 //        (terminated)
		.tx_std_elecidle           (1'b0),                                                                                 //        (terminated)
		.rx_std_signaldetect       (),                                                                                     //        (terminated)
		.rx_10g_coreclkin          (1'b0),                                                                                 //        (terminated)
		.rx_10g_clkout             (),                                                                                     //        (terminated)
		.rx_10g_clk33out           (),                                                                                     //        (terminated)
		.rx_10g_prbs_err_clr       (1'b0),                                                                                 //        (terminated)
		.rx_10g_prbs_done          (),                                                                                     //        (terminated)
		.rx_10g_prbs_err           (),                                                                                     //        (terminated)
		.rx_10g_control            (),                                                                                     //        (terminated)
		.tx_10g_fifo_full          (),                                                                                     //        (terminated)
		.tx_10g_fifo_pfull         (),                                                                                     //        (terminated)
		.tx_10g_fifo_empty         (),                                                                                     //        (terminated)
		.tx_10g_fifo_pempty        (),                                                                                     //        (terminated)
		.tx_10g_fifo_del           (),                                                                                     //        (terminated)
		.tx_10g_fifo_insert        (),                                                                                     //        (terminated)
		.rx_10g_fifo_rd_en         (1'b0),                                                                                 //        (terminated)
		.rx_10g_data_valid         (),                                                                                     //        (terminated)
		.rx_10g_fifo_full          (),                                                                                     //        (terminated)
		.rx_10g_fifo_pfull         (),                                                                                     //        (terminated)
		.rx_10g_fifo_empty         (),                                                                                     //        (terminated)
		.rx_10g_fifo_pempty        (),                                                                                     //        (terminated)
		.rx_10g_fifo_del           (),                                                                                     //        (terminated)
		.rx_10g_fifo_insert        (),                                                                                     //        (terminated)
		.rx_10g_fifo_align_val     (),                                                                                     //        (terminated)
		.rx_10g_fifo_align_clr     (1'b0),                                                                                 //        (terminated)
		.rx_10g_fifo_align_en      (1'b0),                                                                                 //        (terminated)
		.tx_10g_frame              (),                                                                                     //        (terminated)
		.tx_10g_frame_diag_status  (2'b00),                                                                                //        (terminated)
		.tx_10g_frame_burst_en     (1'b0),                                                                                 //        (terminated)
		.rx_10g_frame              (),                                                                                     //        (terminated)
		.rx_10g_frame_lock         (),                                                                                     //        (terminated)
		.rx_10g_frame_mfrm_err     (),                                                                                     //        (terminated)
		.rx_10g_frame_sync_err     (),                                                                                     //        (terminated)
		.rx_10g_frame_skip_ins     (),                                                                                     //        (terminated)
		.rx_10g_frame_pyld_ins     (),                                                                                     //        (terminated)
		.rx_10g_frame_skip_err     (),                                                                                     //        (terminated)
		.rx_10g_frame_diag_err     (),                                                                                     //        (terminated)
		.rx_10g_frame_diag_status  (),                                                                                     //        (terminated)
		.rx_10g_crc32_err          (),                                                                                     //        (terminated)
		.rx_10g_descram_err        (),                                                                                     //        (terminated)
		.rx_10g_blk_lock           (),                                                                                     //        (terminated)
		.rx_10g_blk_sh_err         (),                                                                                     //        (terminated)
		.tx_10g_bitslip            (7'b0000000),                                                                           //        (terminated)
		.rx_10g_bitslip            (1'b0),                                                                                 //        (terminated)
		.rx_10g_highber            (),                                                                                     //        (terminated)
		.rx_10g_highber_clr_cnt    (1'b0),                                                                                 //        (terminated)
		.rx_10g_clr_errblk_count   (1'b0),                                                                                 //        (terminated)
		.rx_cal_busy               ()                                                                                      //        (terminated)
	);

	altera_xcvr_reset_control #(
		.CHANNELS              (1),
		.PLLS                  (1),
		.SYS_CLK_IN_MHZ        (125),
		.SYNCHRONIZE_RESET     (1),
		.REDUCED_SIM_TIME      (1),
		.TX_PLL_ENABLE         (0),
		.T_PLL_POWERDOWN       (1000),
		.SYNCHRONIZE_PLL_RESET (0),
		.TX_ENABLE             (1),
		.TX_PER_CHANNEL        (0),
		.T_TX_ANALOGRESET      (0),
		.T_TX_DIGITALRESET     (20),
		.T_PLL_LOCK_HYST       (0),
		.EN_PLL_CAL_BUSY       (0),
		.RX_ENABLE             (0),
		.RX_PER_CHANNEL        (0),
		.T_RX_ANALOGRESET      (40),
		.T_RX_DIGITALRESET     (4000)
	) xcvr_reset_control_tx (
		.clock              (tx_clock_clk),                                          //           clock.clk
		.reset              (tx_reset_reset),                                        //           reset.reset
		.tx_analogreset     (xcvr_reset_control_tx_tx_analogreset_tx_analogreset),   //  tx_analogreset.tx_analogreset
		.tx_digitalreset    (xcvr_reset_control_tx_tx_digitalreset_tx_digitalreset), // tx_digitalreset.tx_digitalreset
		.tx_ready           (tx_ready_tx_ready),                                     //        tx_ready.tx_ready
		.pll_locked         (xcvr_native_avgz_0_pll_locked_pll_locked),              //      pll_locked.pll_locked
		.pll_select         (pll_select_pll_select),                                 //      pll_select.pll_select
		.tx_cal_busy        (xcvr_native_avgz_0_tx_cal_busy_tx_cal_busy),            //     tx_cal_busy.tx_cal_busy
		.pll_powerdown      (),                                                      //     (terminated)
		.pll_cal_busy       (1'b0),                                                  //     (terminated)
		.tx_manual          (1'b0),                                                  //     (terminated)
		.rx_analogreset     (),                                                      //     (terminated)
		.rx_digitalreset    (),                                                      //     (terminated)
		.rx_ready           (),                                                      //     (terminated)
		.rx_is_lockedtodata (1'b0),                                                  //     (terminated)
		.rx_cal_busy        (1'b0),                                                  //     (terminated)
		.rx_manual          (1'b0),                                                  //     (terminated)
		.tx_digitalreset_or (1'b0),                                                  //     (terminated)
		.rx_digitalreset_or (1'b0)                                                   //     (terminated)
	);

endmodule
