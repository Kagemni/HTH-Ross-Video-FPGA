��/  $�K�=]�Ǡ��N���e��Y�!��ؕS���dR���q=�/������8�|��KۄT=�͛D��!��̍���>Q5-�����k���ͽ.�ޞ��4��&��a匿c�<���)����zu�臶���R��'"8H�\7\�[��jcs@�3<0"I��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n��=d*��O`���ar��x����Y��剰����Q��ǀ��vQ�ށ���q������������0�8ο��6/�E:��3�b��~�;g���G��Ky�zy�cB���q:�cڇ{E�+Td�Z�nF��07�Q��P��	�v�wk��+��Y����`�ǃ���K,�U��.b��p����9��,w��1�⛤��ɺ8� 7C����_��̰�Y��ڭ(v�Li/m�2��eŵ�-�|O�Um��̙��k|�^^#����mK�m�!~��<Q�Wi��m��g0��g|��j��-�.3~E�E�&݂�@�db9��_�2L��}��K�~�����_�ȴ�p���z��o��E`M|���q�t��iLx����t���X@���m��*N^������RP�-M���B�ksl�^�-�2'��Jd杅�,Q�1�4?q��>��������:��op�\L��%�q#cçuʨB��J�;6���d�POS�]Й (X��9������q��!���'[,����/&�:�9l6�Jk�$���Jߛғ}�H&�Ǹ���;"yg�?�"�88$����fj�B�un��:���(Wm2��������3���ڪ�vF��'M{��lI�%	'A[e�Rf��cxݑ��Ȳ� ���]]��v�h��[*�z�1� þԗm����IS�jԔ#�ߒ2ſL�V�������X[{���}��ɻ�BY�Y���1Ų�o����8){�_#��>*Pڤl��}a�.n��W�[�\��(���~�f��ys���W��Rߛ�n[�Y��c�М����4DoTGp��������
�p$�\a�QxWP�b���/F��͍���z<} ����Ź�;^ۓ�2K"P4aRC��C��NJZ��~�����@��M��V��i�&�C���%�jG����p�>v�T��!PU�W��t��0��kFX�e����F/�|��]��w9>8�&�	��(��Npa�"��H0���OD=v��	����Gr�ɦ���ݧ&f��;���!j�����6���~h�7�$�ц���<}u�r�T��7MC��k.���?�����"(_�=$a��@/�$�Y�>5�u�8�2�dVK�� P}��[��r��(�8	~�5�H�Z��n�G�M�>CV�
���7*��צP��mn�K��-Q�(kt"�����XFO(={�"�Ҡ|�E����������%e,|X�<�匌)gFG�>��z^	e�T�Ȉ�g=��|�V�z��U�e+��%i�H�w�{���~t!��li��e
 ����̱���t��ӴܶNR6���I���� ��,�����cSՓt_�Gܓ��3Hű�R;�Ѵj�]��:��,�h@�^0Dي�٘=YV���/4��śQ�a��3����xd���NgM�?<����-v����|;5Ay&�KD���o c|^z,y$>Јw��G����/`?��=C?h���n]e��7��:ݽ� ����w���k��.�a�c� �o���!Gk���L�����h,W2f����e�C-6v%#������/�.u������՝N�hG({̋.�d�)h�(¤�O#֣�B������Y��f�u����]��)�}��i�e���څ0�ߩ���{��CS/aq&����p��D���E�Th�,�s�:�乜�{x߭U�S��:�׾�IQ)��Pp�y�_<�L_�IJ��ݧ9�
^#�Ӑд��K��=�ݎ�̧wBK����t"�웜�e"W�<.-[�	�7���w�C�A��&c1��w�0Y�_�V_�"��vI!�$q�+�C��=�2���σ{H���g�ԭwl���D���N��КE3uQ/^b5Jm!­�^�<����k��ZK�|�-�9A�lv�[�'��*��,.�8+	�6���)�����(v����	�:K;��H�_:p.z$���z�-��rc�b��0Z��f����"�oł��DD(֌����m�P�6l}N����K(��>wL������0H��[���k��2wok�P�������=��� ��1��\KKhSX;m+s�Ğ0GNeO�5�s�ah�)��(֭�4��P�998d��oX�)�v�-���n:�~����
���m.��1|��-a�D�3�PX�7pz��nx)ˇ�N@�D���?}q-X"N�)���gB��69SUS�Q�8�}Q���%�XM��R��q{�H�;f�T���ɕ�'r��t\���+D���z�^��\�C����S�&����U|�B-`i�gK�ׅ��>`��ͳ9�RGe\�B�
}�ګ);�y(�g�_8�qΦ��J(�-K,ȇ����Êp�{��e������>�,e�d��LBjz�V`?�����{��?8n�0̿�:�-�����#���X	���D�' (" ��ZN#�ҫ$h��2,���G�]�f0���O�k�^�?������Z��~�X��9���
�J��u��SA�+	�ǵ��_Nc_���,T�ΊoY��܆ɕR]�5
h�'�-�v�-�K"hh0��S�q�*D�nF�l��go ���$�C,���Hdo&�qh!�d�� ^�S_�۷6aClmKtQ<�i�����",pL���̰�[XzE4Z��~�����=�`W������c�A�?l�nr�3w����|��������'�6Q�fq�w(�.�	���A�4�P���x���z�3�ޟԟ�ׁ��#�[���%4�'���m;v�D��s�5�9a��V*k�Q�`�n8i��Gn���qz�i�@+#�0-��-������&�Sk17����cF)�Q0��"!�m��ms����wS���إL��eaa�}�/nˉ���6��+#,/r'#��sJC��ل<<�T�GA
�;��1 �!ߊ�8�6��_�N�S��yڕpF���+��nP��
�A�J�UC���l����'"<TH�� )4,��<��"FD��=%B@���py�7I�"��U�oei	��w�c�Ō�`sX��������ހM��5��4+R!�\�B�@��K]����^G��®~�w���Jp�2��UZ\��%��V�"~r��ڗ�Y�`h�3 e�da������Q�m�,��W���ݞI�5$[=�л.^���#�I[��_�{%�Z(�f�c�Pt7Z�pgI9���P ��$�0K�-���#�ۼ�̜�����5<4˒�p���K)r���rXcl���9\,z�t*�Cdm��-p7��̑��2��*sy"��ہh>��F�+pHP^g�����f�C)^��x���[M
!��I�kj�3�UQA4=2*kN�~}J~�orҨ<�1������7@�^Gm�'\�=���C�J�/D�L9�>u5�7���s?)=I����<���~�'c�;ن�p�}(��g����td�����;2���>�-����hF��tʁ��U������g�_�-#�1����B��h,��?q��8�C������H>��z���y�s��8��X��׭g¥y��zߒ㰌��Un����]%�F�1�D,T�豠G��]A�J8�=�)�A�����zOQ��֧�ZhI�ҏ"ߝL3�&��Z�؉ ��S�4���L��؉�o��{���l3�����<�]}�D���z`K�b���R<(����a1ޫ}�ة���A���`����|��<8�.�kq��:X �W:l?�<r�A�W*k�ح���_��׼���j�}=5m9-	�pcկ��i�nf��2%�	���o��!H�ψ��7��
�%3���)��h�51=�x��<XZ�}a��O���vC���9���@OЗ���;u0V�8G�M�F�"��xOpؠ��GHԌk ֖
�+��}�����B��W �<�����z�gO�'N�n5�S�{a���RŪyi�F��nZLm�<��{v[�"�15[/�+&��)�˱B��GZ�O��%�$�d�^-��ދ���������Y�xЭYj
�~S�U�=�?r�)��`�r7<�T��\�_o�����3�4 ���2̈́x�k�v(Xo�$�UG��)�r3S�W��o�논'|D��2A�#��!��5)'����]Qճp�-jɗYÝ}��Kg�)����"t��a�0%�m8�竘:DM�����;�p*	��Oh0�hE�1�9D�D8 ��v@��W�ǿJ�a���%E��O���tZ�*�����A��t>���gX�I�:����VB��o(@9g�B[p%�G�I�EX�1]�DO��QzW�j"v�Kɟ�v��]�y����k�g.Zo�n�:�/R(q�uK�ж@1<k�	o��	�;�{�yJ�><h(�a,=[LQ�E�M�����t%n��x\��$X���mfc� E�L�:9%�'e1�mrm�ա����TeM�D�x���@U��n�	�3��� VKz�r��1��6~�L���RQ���?�^"&_���G��ʃQ�rb�-!�R626�3��S�f��~�8&������"yL�=�p4���
-��c����y�IIy�G�#�1+r�h�d8�U�xS�����˔}�j�윱ܟZ�B1�E�I�e���_b��Â̽t�
��H�e�!%I��`_?\#�b���{\fq���p�,f��|(�0M����W�$^ђ�ɇ�P� c�P�ę�@�Y�V�5���)���f��G��Xtn�Q����HC��yT�*@8�Cy��Q���]8ҳF[nk�88�zڽAm��7��D�T�PQ���l,L���7�a�6����:CqvB����N�ڐg��$֟9������D�� �ɚ�?�9����d�S-'��?�$��7{�"��+ek��:`�I�n�Y&2vh�݇��>�}D�7�#�����dt��^���	9��1.�௓9b\Z���tϘF�*��#F�+��'d-�+U*��0Y��o��y�֩`p�͐��%����a�t�6N���4=�D�?��%5}e�߁Y�)Io��W�]��H��@�Rr���1�9��a�{�kpw+���K],u`P���4�z�e�K�$�����1$�(��Ƶ]��9�KCA�!�c2�.�`���CC�7b�t����i+}|8�h6��\�GM7��o���4a��ߡ�ϟ�����v�|��A��g-.�rT2ŜOp�Z��6`������䤕���Z��!z�d�f�f�Ӕzdf�!�DWL�-���c��s������d��#�D-{�0O<�6|!O4*S��?�hf��M�hG��lG{k�Ϻ�j�nS?��-��d�>,��xk��f��[r=�_l���`!r��	P�>�c8�+2>��lEP�N:L�d�QC�^��[e�)Ǹ_�/7�V�HD��%��xsg)�����vB��>�mS�)d9L�\d!ZW/��^>DY&qS�@����QQ�Bᎆ�v.�b�9s=g��b�^ִ�U6�Э�"���4��B��.�_�/�F��ɵbO� 8g���j�o�����@5�Ŵ0� �9�n~�����7lI��!lk�O�
������*!/����\b���/g�Q���Cl�9b�TZE�-�K}��Ȋ�w�V�F�:M�����@Y�@���b���D�BSP:�>��M��[�0�q��pFP �aEg�JS
�G+}ͩ|��ٿRM��j��	p˗.�*����+��{����$
si���&�r�������s�4�T�GiTO8���u���k�����1`��V�^KܐM��]�_96J~�}A�����zr�W�|����$*�-�)���ǣ��/�v0��}���/��q���|�q�_5�*")d�1kй��%�\���7*�#Fl5�d���p����8Q	w���l��#�Q�Z��lf�vn�����@|���!dT[����ҝ *� :��sϲ�ֻ#���wyw$Q������&�,�D��B��^�H���1!:�U��zM��V`;;q)�k��Khޫx99t�d0��y����ii(u���������7z�A�}�G얯��kfˠ�I�n�/pOL#p~a�R;g��ԑ��)a X�#�z-W�H������ҼZ�ki�y�X���У��
������V�9�G_�[����kW��r�ws��nɰ���ZHOI���.�ᙫV*��s�8S�4#$ׁAx���얏����g˰v��~�*U�.{������<���d�����ҁ�#�uq�8��-�����O�P|�����wd,���]�9���h�����p���.��c��o*������FŪW��5��B�L�:^g�d��cr~!�/���[!SKׇ?
(��L��Vp�~zS�0+\v���-��<���a�Ce�?ܑ�CM!]>2���m��g{�oW��8��ro)v�EA8�@�9��|�z������q��=�^����߀�ӑ<X�Iٵ��E���i#��.tU<��Q����{�0�:_{�����V�l����o���=Mj��lO:ļ��-n��[���^B#!����<�`�+��2�aH]�z>���"\�C3�.rYS|��.b�\�!u���ay�k����V͛5�_I�4��ׯ�C5��:��s��L=9B� �d�m%Ş�D����?�F4]��|u�OR��*�UO)��m��F'�t�ᛋΓ�D���mh�w��lͽ��s/4�� �r7Q���G�>�ʩ��wv[Ugu\uT����Rؕe���n�f�J�l/|�+G�sA��F�|�e��r�u��{JP��k���\�İu;��y;n�GAWq��Ɛ5Z�#F����#Qn��:��؛ s��i}é�ߠ?�(�6���ib+FB	[�:@����������᤯1֐%�,��;��r��bU�*���� ��8�@H�g���I�Q���SV:���#��D�c�;^:D�]L)��سzS>*�ɚ^{�8���*��
i �XeJ�ɷ0
�z���<�b�Nޤq���b�v��ҥ�ܬ�`���f�>i�z��4f���Q�%�W��D$��ƞ>�&!)�r�}��^��ℷ����ed��o1(v�!_�}"�w�8��W6�3K6�q⺿0i�J�#LI1�KϱSc Pn���=���B�i2�(�n�U |e�������%��.y��}Ң5���p˞[m����R\�������8�S�"eH�|�����+����$�4��\�X��J�n'9�� ��٩�7WYe�� 6g�.��TK��XD���P���C%�7�uO��&�D:�]����p�\ T�3#�a��h�G����R�]�7�d�c��D�=�'Z�㸒?S�[��L��Z�9�̼Q���("v��	x� �u�乳U���s¾���tA�������`ڬ �G"�Ojb��2 q�q�!\c���nK`S�`D��l1A ���'79P(����w~�v�ДќX��ֱ}�f�I��P�`u����oz�:!��Y�
����m9��"�Y�'�s��)��O(_�T�E�U]���������v�Wc�yȑ�	�l�&�!`ʼ�rL@���ZC�qd�K�y��y\�G
f�z9ט4�ZZ�4�^��I} F�.��,��� um�"�n�	k����&4�sM�l��b�Z�����='VK44���=#ژ?��-N�ͣ����ub�k+x�f�u����p�_t�U#�-����"�4�\�L����wx)��Pa)�����������0�4t���tq�;��I�Y~���h�K	�c��ŀ�q�7"�ԯA��e�{͌>��`�9��M�����'�W������jK-� 'T-�`Y��;�yH��4��ce�~'�aZ},����E��n�ZGL�O���u%��1�� �qV�1?B�mn���܌	Q�L���ꪺ�S�1�+�2�E:�܂��`��W[��򷞹��!ebq+�����\�����$�t��&�ͫ����ޥ���O���F̖� 5
�P�LƏ�oBL�\�E�{iWC�_����^����1�4Շp�
�8>��X5�����#�!k\=�s��y��s'���@����ll&�|�Ǧ��VP�G����B�k�2�2<n[�1=#����i��>�{R�13~�t`�U�����[ʻV�0�DA�p)�l�Nw1&m�vJ�n�t?)�v����lm�U���ʮn����/bh���G��MJz����(q�TD�/�q���h��-|�pC����w�XC����΅��tc�p��0���G�䒾6�����7a"4�G����4����¤s��y/D����n,{��桐7Ci9���gp��������$�:c�zm�!8�B�pS��jg��;�A���`�� �|�3.FK�}ܘc@�.��m^9�����b�pyDL#�`P������1>C�Ò�!�&gz�8K���3���zUA�!����� ������@~���;�5O�U���'��q8�.�:U��X��ĸ'j���Ƶ��oj�-=^ !�M��1{YP>���SG%�c�L���U�7�پ1_H;N��Ȉ}/�p�4KM��r]��/j���ݘ̓�g�+w�����i��#��;>���Z��!��(���c/?�.o�(�넚��rr���y���&��� �}ՋB��)��'P��2]��K+}��Y��N��*���T%��Υ1�}��F���ePzn(�%@[�v}L��C�"�Q�q��/]�.��f:@�08)1Y�<Ψ����Qt����;��0�4PF_g|]�8��gds2��K&��B�Y�E`V�e����I�JG����Q(`�N�~Vq��.|ٮ�XwZ�(v����c#�o��5�6Sb��A�G��$����T���Yk���Ǉ�'�a�<�����#����J���܎Z�!o=�t�����ky9�p%��R�{3�#p�M��z�Aw*?�Q��
�rcH)`����Y�D�`�"ЩV����.�|\�(�]Ҡ�����ᄜ�;q'T��:�u8>�pd�},J}�.z�o�;>����:�J;#q1���S����.*�����(I����6+pNf���H���S9Ӵ{����%t$3�ÆE��~��Vz�3��m}jA\p�e��n�>���s8��)�4�g	46��LK��{Ǚ����r�Yt�R�a�0�'�0�%P�ɑ�_��KKjh�������E��]b1�p���SY3D�
��d�tBu��hy���I��`q!�NA=��/NФ1U(h��Th1�x8p�|�F�)�%����eը>q��^�m�cݣ���<��'I�ye��c��d���v{�x�����*��w��At������-�_�g�EPa#ߴ�����&�}�#GF�!�7�'7��,F|��G����&������>
���s��P͏��	5�ܧF�]��h5o�.�P6jMӾ�}v[�2���Qmۓ���3(���f�W���K�.�qRԃ��j�a��1��-�`˖���,2�
��o��Y�43���f��e���v
8���u�0�r.�J)�AV�v���S *9m��mN��D*���D� $�|��"�QX~���ǔ�+~`]��L��J�9�hGw�0����I_v��'<Q/	�M��ܡ-6�z���T� D�6���z	Y�y��#�ʅ�Pw�5�M�*e�_v1�a���h	n��!K����\�_��R�b�5>_(XgV��μ�����P��U����$�ēR����)��}Ve�����$�0j���a�����\�f��ٿP���fc��lȺ�#��ɥE��9GCl�7X�fzM��H��{:;ː�&�V��: EGwiJ35�n��YIûp#Q'��ӷbF恟n�i;9��KN�ᾲ��-Kv�r���&ljMhuX/G$P��J͢�ҶS�� ��Xb�h�%��x��<�T�˩� @��k�۾�L��� �(�_�0���+���������zG�\H5����:<����l�#�t��`�����P��|���<���<�ŮK`.���럙���[u�k+��y�A�2���jA���%�TH ����K���Az=��k�$3H�z���L�a�_�۸.y��r)����fU�v�\Y���4m��>����A`T��C0W<�+@
���,�,~���v�JH�AmP�*R���<o2�zS^Ӑ������EG�Q����5�+�>����>��=��](�k�hj��Ĥ����V��5-�R@�c�G��0�C������l�������ZO�o�v	KKO wd���I.���+B=#��p�̽���4�H�����4"N@i+ܷ��	Dc1@��H<*���"��X����-@�%5�u�Z�KV�6�/�� �tx��n엑�F��\����/��7�R�'��y���������*|=4�����&�\v�3T��5�rW{�.�C��2a�0�