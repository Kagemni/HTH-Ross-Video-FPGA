��/  m�u��\b�\�:a:�#8iAZ�!�Å�g=t7��_a��&�cl ���
�#�J��l�,�\�1��'B���X��8��NH��������ӎ�	�s�
�#~U�S���	o5?��P��4!6��O��.F��r}+��UW5��),+רD���nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n�W��ߌN��5=�8�:N|���gp�P�ظ��U��)�& g�J����[��kC���Rm�߽F��oot"��QM_������,r�� ,ǆ�{E#~L&�80QMa��avXa�*_1��@Y�- "I��Oh�:�-�}g�Q<�����]v�$�:G�#��t�����j�w�gtGGK���K���K8Ù�@�F�~��7���㕹�â�N�l���&�ڍ������ME 3�;%�5S���{H�d�J��r	�cH��g��ͷ:�3�{>�)�u��+.��ؙD��d5�J��P����qS(���p*dB����s��'�.ޭ�����۔E���R����`��](m��ש�0)P�K��Sϡ�u{n,��@X�,�s�\~S3G
����y�Ր%�5�7F��s��\��#'l��������n��%��%T�P]F�UF��ݓG��O3�/�[����N��o�C����������"�d�w��u�(rD)����W+�	��8�|\S�+��+�	���,/�M�vo1f{����b@�1�O��Y��֗�6�i��x���6�������V�"fy�Df>ڳ��K|RF���Jl�G�r*���
RǆLI���UY#�"i�
�7t�'���f�#T��
�/۫���ќ�˼>�,��o�_����������L��2��Y\��Š���j;� 0)m��Bh�~�:�a(��2վW׾�m�;�� �x��қ(A�{��,�U�R�i�oq�D��� #�<&��+���A�����"g����rQ�,TBJ�$]Z35�<g|r��;eS�r�p�o�eH:�2����:w5����e�@8x�IQ���".4I����ߨ�]�9�3m:]Ɔ���<>�̂�=�F-�.�UC��|wD���e (��`�̒����+����hF8�r��t�fɐ}x?�L�F���g�V�Zy M�.����Wq�����'6������Ը���n�A3'��j���ߪ����̸O V���K���&��9[�B+�+f�^�b��XIU���I�g�A,�[�܂;>}�Z����� TC6([#<aZ�
؍���N�q�����n���{b��$��1��RG���	$�v`��P77��#�X�ً�|��x9CqO�N�������e����7g�ۖ�voy���L�� D��`��q.��fA�F:v��F�/)���K)��s���'{mJY-��
�_��~z���0�r��Rݷ�*͖	��0P�|�#�G��g�\�L��#l�j��,iW<�����K����0�j��%сWkd�Z`;x��+�4�NXyU��������LlX<�v�P�V���ji_�V�BG.���u�
� �A	�d�i��J�����߽D�G�9�P���ck臿.�g4�^���OA���޽|8Z��:],L�SˊLĞL��ʷu;�X�Ac�4�N,��fk4U��m��d
u��G�4J��F��(����YW�'2V֡81���o��EyH��$��P빔�.9���@��/�^��09r �����½z�E,����5&ӤB�	�-���ӕ������bx�+N���u��	f���?�F�'ތꘟ��E���,j�в�],	�c����{i��kd�[Ҍ�WpX]�+���6�7L��H]IT��oݎ��I+2)@�u�x]�U��17��B����$�T^Ri��e�$%���v�xҍ��誊�C~3��5�Y�����.3͎1�Ί`S�q�Ȋ���ꓺN�o�ra�F�Wt�%�u���= �&5�.p�"�8 ��WM:$��̷$�W�P	'~��,�h��H%P�>J,5���Q��+ܨ���+���Vn.:��E��q��G��� �:e�$�Z��Y@��l�W��:���<� ��$���x�ϝq}E�0����[�r�'�V0(�i�vu"�v� ���(O#�pv쓃�p7L�t�;z����<�w��p�C�;��Bo���n�.ߐ��Px��_s�Y�e:���8C�S5,�v������Nj��^v���S�;i�����+��I�,�8qx����,���YSu<&���qq�k�,��j芲z�Q9�m)�?)�� �0�k�w��V�W��t���3���ƿ	��Q��?F�;��)-�g��6�P���0�R���wTC`O� HX����;�����/ܞ�k�U��Hv��=<�.�m%{47���GtXH��m��i3�!؋�ӻ$ɫ�z����*�n��8s�ؾ�'#iVZ��?`�+��K��F�����a����D��grW,�H��w�7��7b�だ+�eh��4��!��/�+Yf/�D��WƮ��}�-����t���T� ������-��J��1��ڌy�)@�,f%1|�����ȡ���c��Y�����R6�F�.���<x�b�bh&n\��d���Y��A�Sr��<�A���lĬeY�3 ���q�璺/e��fl#�����������	T�����f����맺������e�ԩ���S�iQ�|&lX(��&mR�,7K.���������|����6�P�����"����^�{G��cX�zܿ�İ���Q��+�5�@*\x/0,�`���dj���Ƚp�����C�~Ӥ���Kz��PDH.8��>'��ۨ%d����jK!Ё��t�\�������Z qεho��:�o�������aop��݅�-���O���yO�{P欣oV(5�˿{M9g��L���c��e�K���D��e!0wNF�9���U�"��ogk�wk������-]�KŕB+����P����G+�S��x.�C�!�)�c>N��%>�[G�\�$�E�ʜʯ�Y�:�c�%?0�_4	���E[���C��,X�<�K�L^���>�e@�Ny������[Ԝ���|�Si�g�!D�[!W2���
v��:��8o�J���
Z�԰�%��o�¹�0�o�ô�`���N�slX�٘_�㱝��Y|ɼU�l^cf����d;C����4A��}u���i����v�����X����	g<~���.�����+���o�c'����	[���&G�_�A���yu�	M�/tm"rX꟢��e%B�*QY��cĖ��������E}��fzv��<�ba��m���I��Ԓ�&I�V�Ov��T����ZћPvE��b>ɧ���1ҧD�������_GB�l�x��qV�US���4�_�	��i����	�9Y`�ဲ�<� 7>&Z��������m>��\�N5�hV*�+$��S>�����*����[�ҧr��1c�,�(�F��ˆ# �V�HxH�i�o��'9�3�qљ9�l�Q̶Ӣ��f]�g6���ڃ���0���b[�����^�,���Ա�����\�?��FK�M��'�e.�-H̕
��KYJ���H��,����k�.[x?S_���ʎ�D�}� 