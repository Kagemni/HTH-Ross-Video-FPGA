// clk125_pll.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module clk125_pll (
		output wire  locked_export, //  locked.export
		output wire  outclk0_clk,   // outclk0.clk
		output wire  outclk1_clk,   // outclk1.clk
		output wire  outclk2_clk,   // outclk2.clk
		output wire  outclk3_clk,   // outclk3.clk
		input  wire  refclk_clk,    //  refclk.clk
		input  wire  reset_reset    //   reset.reset
	);

	clk125_pll_pll_0 pll_0 (
		.refclk   (refclk_clk),    //  refclk.clk
		.rst      (reset_reset),   //   reset.reset
		.outclk_0 (outclk0_clk),   // outclk0.clk
		.outclk_1 (outclk1_clk),   // outclk1.clk
		.outclk_2 (outclk2_clk),   // outclk2.clk
		.outclk_3 (outclk3_clk),   // outclk3.clk
		.locked   (locked_export)  //  locked.export
	);

endmodule
