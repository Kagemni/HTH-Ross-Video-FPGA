��/  ��]I��'|$���
�8l�Do��_ƾ�8�H�a��n�K�U�Ãtݪr��L�,���|Hlr��J�륜'��#7��:,�pj(��#����!��@J��s��3�TӮ��`x����eE�R�p�AjU=V�D�����=���0������nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�UtK��^�)A���Q���=�.m[�F|��]C�9o���m����T��i���`3��.uFh!%�S)|cph$��ڞكRy�n9��;W���|�b
���06�^��'��XO�Y�z�+��^�`R���[�^i��.#.�Hu�!�^<�Z��{�I��1�Ꙫ�r�R�9�����<�,���W��%�jٗ*MG���V��4K�Ӓ}�m �ө���;JԂ7Ŵ*�u���Ɉ��+D�A�<%ZTq"�G��{�RJ�~�ɳqo�EsG��%�;�	����o^.$�4= �7_ka7�h�P�0.=Q�M��T�x�ZG�G��R��������<�̮Ϙ���.�Ӕs	M_�>�=�,�]y��fi�ݣ.���!�}3hV���*~�8Q!v��w�
�QI��1k�Q�
�����y��,�o�yG!D��c�N�'����f�|N��L=�� ��8�meO�[�z1�h��#TMd�\hT��9L��N\�*Ӟ�a�k7�&	#F�Xyԣ�^J�R��4���1��VVw��3��oܣ%��L�7��4��WiΜA<�.�҅ua�c~|�¡,��_P^���f��)��|��$�bQr�� ��1ex�a�ژ~��C��~K��Z̝؃�Ve�o�Bs���I�5�3Zq�1���Hg���)��-W�{^U��wc�t�4�x�ͲU�pzJ֡E� a0���~sM��b1~�Y���Q��_|P��%}s�R�A��wȀh80(-py������X�}d`=�Y�1�G���#���
��h���w�Af>�{xJ;a�0���?MX-�H�{�E�a���j�4�ѭf�-n��/�	�L%W�=&�-���^[�L��+>L&Η݈mNXɖ䘠Je8�Y� ���DC���y�g�yж~�Xq,�y�6%��b{����NKfW�ҿ���{"*&Qm�<L��s!���35s�P��^�)�-�ꥷ��蛗�W�>2׬�K�V:�A��'�HK�z�P�J���w��7N�:+�~�28�aJ��-B�l��,Q�|G�U��M�v�����T�Z�
,51X�ƪ�R�4L��X��y�S� ���CUj�N=M�U�g1��
��G(k��m���q�IS����ï�%���>%�CKo8�QO�*�m�ځ��!}�1��Òq�	�Cdb�I�I�Q��E��� �����ĝ�A��_-Ck釾kd���<��0�C�*��\
9���c0k#r���r1�/�^,I���D�)���c�T����w�c�a�F����r~�m�1�޿�oV"|X�n�捭���ckت��3�9��|���
g�ꆞ�~�����kF�ӝ�R�:L}-"n���!|�.���Mj�<�s�s]v��WA�F�&�T��ۭ�p�B��(��Yde��|<ޞ���Sb�����w s�p���ʇ�<,�Aʭ�~��K�*ۮݴYB��(eT���^��bz%����>A��D�<vP/P�8	��r��$�3eO��#6Q
��6���%�_�_ͽү!��xn�ū��~Q�=&޸,�0���#gk^j�[?����_2|�EF�F��]���d���f��XG�qW��Ư��-[I%���K�W�Z���M=�z�J"J�W�(Wu��;PŠ����0eN)�i1�7�b/s�,���jø���f�N���)����'�)�}���/ΤZ7R�7]��z������]�ٴ���DOA��k�V�Չ�dQ�?�Hd�H��,>�����:�ܺrN���hD*�W3��΢+�㶆�;�@֘!��Y2[';IL�C7�0��*p퓾r����V�6ԱR����w��/��n���s�Ž�?�S'T7��i�6�?�G��`w��
^X�v8!,.�s�>y�P�-M��op��]�{_bGF; �8+�e�2���� �kf3�p��H�L ��2�:b`qx$�j�\��i��
a������kW��_�|�L����d�� ?G�D�#���A0g�_��#��1T�es�U���u:����:p�xF��{�_�e̜]���s����9�9�*�&��}3��]
 �Q"^G��,=�"�ΐ�j��~񴢋<�~0!fa�pm�������4<�*���I�M���co�ө2ڌ�XqyH�z�J�Ȯ[sّCT���Cq�1�HQ!rӻU����&ÀX�Ǚ�JO�=�ƪ(�dC4�܄���/ ГG�8�7��i�21z�����j�n#v��ܛ�a�u��a���߷���m6�� <�$ϵbs_>W��.�����W�$�8�t���h\��$熭Ex��0���W?k�s�̢^��yf��zM�X��b�k�ʳv�!���[�2H��������<?p�c�\]ʱ�o�7� 6*�Ufc��^H�@�j��| �)�=��X�X��ն�~n�{��g�%��
A����9�*@	���2��M��G�Jx���u�S i�������F��Ҏ������O�(ڕ�U���̄�V&��H�k�UH�v��Jac0:�d=�"�y\5Kg-�M�*Nc�D�Hr����-����d�5�E�R|��֑�ظYR%.nId��+�
Nn�,�WJ2�X�C��jPN�a.��5sM����v�7�����j6���5i��)�30���t�k�->t�����y��+�&�N��0�Ws���(`4��gw�f W�p��4r�c��tj)��Z����*i^Q�ceC�U�De8����R5�W�l;o�OM�ʔ�_�;X!i�p�{���+��k��0�9�=ƞ�������QāX�=4C�D�a4�\\iZT�7�q�7�p��2_�@=�9�q�G�aluz�[;\��y2Q܂Ϙ�T�H��&+�mm�|�{�JĞ�	��w�k3��k�-�iF���#Pg�� ���NGp^5[_W�?ٔ��DƐz�_���3�����&`@������ ࡢ=?^���Q�D;\E��e��bʪL�<�Y|vĠ�l"sR|�1$�u2AP�����v�_��<����t�K�w���mD.i�pW6!!��la��j�̢����¡��I5�@#��d`�^nG�1��t������y߱��a���KM�(�xF����O��M�%-��Q�'	�8?<�W�1 =��x�$�RV�8��i+Ƹ�*�'y��P��:���A�c:�B���1���G�(��21��|j'�!�=I���S���SWAJ����тW�vrХt����А��}`(�ꁬ�-���3���f��H��h�pW��Stg+��� �(�R(*��7�V�N������d�l:<l�1���8��R��J[����U3��m�dN�Xo�d�#H~�_3�
����3����>��X��`�9"��y�C'����.G��s�U�^0������$ԓ4D��h&$L;��7�(K�,�մ�1��$
�r���8��qG��n��L%�3Y�c�e�c�*��3%��E��̂
�N�m��^-��L�5�;�1''�K�l޼�|S����ǒQ���~�;\\�4����N��m�]�������^����\>x�[N?F/:[��#'!r��M�Wՙ�b|�g�=<0�_!�9�!y&���Hw����u��خ�R�2D���w3B���|�>4�@�nVӼ6|����U!� �D�՗�Lh7|��D2�K!<h�o�̭�-�Kzi���A �R�#TDCfzN�;CNEi��+h�\zQ���#����7|l@q��٦U������b�gT3�q��Z�٨�G/4t�q
G"F���M���*H��hxRQP�[{e�:��� �u<�K�����o/�J�Wg��Z�q#��d~my�I� ���d���Du����~�'}�k�G�y�ia�' ������6G�E<!��Ӆ�d��Z*��_�j@����� o�6��F��#��e���xӑȶ���և��Qx�|�|w��N3�P�V�|;�+l$��q�8�k��_[�cd�E��)kS�*= ��>.�αT��{�K_!��xa�`P&��Kʡ?�ɲ��G��o�3�f��	<��&��d�7�C[r���m<+Cc���pZ�&�-��1�P����%5��3K��B4����ڥ0*?|�K���E��	r!ä�ŭ[���Q3t�*ҖQ���X��*t	x4�z�F<ߵ��z��-Y^�["6Y�׎XJ_f�PN�%�=��L'�;�$d	_Mq�T��N�V�dG1�M��L�߅XC�}QݽL�b獵�(Rĸ8� >��o�{�N����dgFn�:��ݓ���{�+4.ݵ�رc����Fؘ4�DS��hHP�\z:�ey�� h7�b�$G@ ����K�>D����6߄Vhus	�nR8rA��N��x��V`)7$�Y3
����P�-śBw���(*�
�e�wZJ�wߦ*���lWԙ޲��=�����93��~O��xI����ܐ�D'�	�7�j,�g���KZ��:��Ĭs�;o��u&�1=�)������Ϻ/�]7��S8K��t���;�{��'����k���*��UX?�㪖��b\�� �f��2�'����ɰX�arN��Q�avAGhj,�Z6�*��P�lv`���g��&�7ȭV�4Fp�հ.T��Ȯ��Ɗ:d�1o�1��i���ލ[��N�kD����ȕ#��qԷT�Ҕ�h��pڴ����h;,mfc�TC�������@GIl&�7���E5�"�d��d�e���-{\՟K� �!m�۲��H���S�u�#����.�c�_Usv��-h%F��ܡT#��4�3�]��*������T8yK(��y�qB�X{��o�m����EU��BFf�+����@ Ÿ���ܖ��A�b��^/`����M��g���þK��W⤦_�Kp������{����˿��3
��o�������q�	���i��r�%<9!�PW���U���!�c�D��1�LhIÈl*��Y��n�Oc�Y�3։K�o& :�;�>)(�Z^i�:<�'���	�,p�Q�S,5t��^��-�/W^��&�Ξ�����2�iҌ?A�j��|	���+-�.��m(�~t Nq0�/���Ԏ�)�_53_y���<H6��	��Ŝ����nNce�F�uȨ ߟ��b�&���3ʋDrB�R�p�6�P0���;�`�J���(���ȸG�yy{�փ�z1�r �°�������(��Y��bNژ���.ߋ�am�K%'�~�6N�Lw&P�d��+��ry�g�"Klj��%���X���^�3m8k�9(!uo~§С��V�)"Z�w>Y(8�����`���o�H�J���i����K�R��N�����#�B��`�]WN�j�۲�C����h�8EVd��o��`���(tg?�Xҹ���O5&?�]Y�|�|݋|�C�7����>�����d�%�N��mi!��Ctu<����e�����.HW������m�v�'D��]�	g5�Ta�OP)�a����}�Ax�K.
�I��\�=v�s�u�u����f��H��BOU;H�>�p�ymp���{0�5����/�4�G��ܰ5�hw�Z݀!x�D���aC�I�0an�@N����Xhʙ��]� @�"�<�L���Z��	�k<q?�������V��g{ �θ:�ZF��U�$��l�g�`�\��-��3�K�e�9�`n��5�@���6�1|�L6m�|^�� �!-����G/r����yOF!�)���?Y"u�d�h�<��奻��	3	9�퀥��
�x��9V�[�������gG�������h�+Yv���E���/�h�f��--�n�W�m/�y�~-7�Y�H���t��6y�!��^!×T:A�4���P�~q����t�7D�&36q�������Y'���h$/�1RU����I�6q��D�S��ɕ^����l�@�����Ӳi�)�����t�
.e���Zx��,��J�����w���[�����g�e+������B�"�$y}��PY6���/�:*#L�z>��$'"����Tr�G��1yW�5�2�ZU�^��߬��g;i��'s5���T*V�cˬ�L���B����Y�A�cJu�����R[��� 4N@��lY&Ҭj���.PI���0��D�d(�iuh*��h�Z=��:�yt�i�y��P�ֆas�s�8�Tt�ń��D�A0/�4���z��N��>dF!�e1��b�Wp�4��;?�U�J�&t�=���?[�I�*fi����R�'J�T]�����Z�gk�#��'iKҍKi��4_I���Ab��ƀ��ˡ^�p�NOy/X�~���J
��}��Te|"!Lm! ��LU�ꭤɄp��́Mj��a�ќ�H��pqmkr���3���$f��*N��r�vR��� h�d{3^
��v� 4I�Ic3��?�G��^�(����ì����Ur`�9@���7a�ߞ��L����7IY2`�16����?#�+ ��@ �ʝ��䖿����ls17����Mݥ��&��_cmC�*���f�jֳ6�g*�պׁ��P�CcEN�d��ԸI�Մ\g�R�ZF�)�1BD�4�[+�6˨���1����Z�4��TGE��٨2DC���`�-�T�M,�Cط��xN��TFbD���{��Gݨ��܁kgt+O�5q�L�{l-=�``ߢ1��O}�(� ]ciUx}
d�CsZy��zh2����k�2�1M���բ�8R�vq���6���u�����������eΡ�͵qM���P3`�e's����l, � w�ux�pV��f��,��qť��#\ljӯ��N�u�c[�Y��̉!cnpx�ł����$��5��ҕ�lO"�{���2�@�N�����#B�ء|c&��<����u�(y#l�YX.濥7�����1��;��m�w��>}?F:���mN7m��pQ̘)���,B���$�,�2��u�K��P���X�	Y�U�Ws�)^��7�F�l�$�2����s���f��jX�,Z���z�����E凨�+ar��d��׼�Ra��M�,R��!�RrC��JG%q��ZC�"�f�Z-�GG�Rsg�wE½��l-�Q��W���e͏�9v3�gOm�7Q�ʻH�x����X�u�Cf~z��bЅ"-T5sK�+��?��C6��x"�0#��%��J-:L��H_6� �	��l�s§q���Y�!�<9j����ȫ瑔Kt
8D[��8���h��x�	t%��G���?�����-��o~�84"#t��h{;�ʌ����<�ʯj~�?�R
?�#��K҆(�k%�4Xx�S-F�h�j^�0<�"S�|y��(*S��/��qPap��:�qMy����c���`z�O�\KPd��C<uĮĭ��,[�zG�O�A�
ZQɞ�6�Ye4 �@��-��Ls�tW�?\i�9~�Ĉ�:'2�$��֡�~����%���2g�'�(��q/�I��Y1��!��K=5�\1���q�а�����(��O3�%�ʚHϣf̚{l����J���\��]}��1i#�~�����u5e^�@H��:FSP3x��ńo�a�� rrz����T�+pf?g���p����@��ā��͂�{�4�{�_�?m�b�/�1g��g�ňj����\+-�u�1��f���&����h������>3�%v)���O���N�u��픁l���SlV��|�P�㿺zo>�F��M���;��J�W�� N��ޖt��8��S��/L��O�caL���3x�e�Ԓ7�UQ!;� ��\�^��7��X�/�����PcuB�����4�����^�(�'��p�c���"�0�Q�T�х��2 �Eܕ�bX�Ȣy��F����`�m�>�����:�)(��$����/�=���J)$K����: �Z�F��ޛ��@�둻t��H�X���� ��ƛW@�������� �_BU�bD�W�w����,'�T/:i٧4�9���������u*�!-����F�6�5��/H@�L�5�1Q	c���̤O�! �0�pպ���r��3�v#&��ȞW�xtg���`�1�k���z��t�V%�����{F�2Z~iio��Z(�O�e�}f��H�3wC�#�*�P�A,B��jy&��O�C�Ю��{�1��PD5����{Օ�A����E0�xeLM� [ҾF��-?/zol1+ݱ�l�8p(�t��<ѽM��i�@�01�H�vϠ*�8��t@�����q���KH�\=�*_|��G��r򚮭LTP�F�=^�4�(̍��JQ� 1"�'�qh[G�{�Z�5X��~�(���ű��l�Vs�]y������O.�w�
?�bE��`���7���ڟҞ�l�7p�d�8��U;B���C���#�ps���E0_�H�(���oTo���9�H�^4Yrn7�;��ʘL�p�i+�u/I7ljm����ݽ�չ?`��7$h�4��ɮ;qh�h��8��;KZm���WW��i����q+��]�6B"*-�Oҡ��u7�r71U�4A�����Q(3�E������x��N`��xD�ӵ[�a�n�M�C�՜Z"2r|]���;�4��<��Tw���A#���
��X�qMw!�ъ���񝫋6���+b�?��+���ʢKmQ�]y���.ɓn�s��kN~,K�;c���t�3BO���.������^�y��)��ګy`}���v�^0q}&r�s=�x�Ym�-GZ�e}N,��/,����`�N۫*��W��"��w.��E��A����r�}��e/��:�f����������U�:֯#�{Ck�Y�TH�ݶ�C��6��;�� Pl�oin ;���U���u��@8&�A/3۪P9��_#��Gb�S{�=�����j��)�
�pE�W�^��6ɿ��^�G��B�Ȓ ����`���� ���#����hl��Ifw�{���\K���t˜��-b�%E)$����T���=�E��*.�XKh���s�-~d��f=Gғ���n��f9�1+f�C��u;�[���鮞M'�5YC{%��ީ�t�+��಻���L�ԕC��C�����-�.��t�G�����r�N�aQ6�U����XnQb�uH�)@�E��;�z�b�S���@�i*���ĭM�����E��.���:�ݫ��B�1���no��y��ZZ��TL��A�9�8�%)e�|K��`w'?^]~���Q@�g��w3~�0�tM.�	q��Zt�)���7�@a�r�Td�� ���s-zl�|ׇ`���)�Q���s�`�7�u�?�=0�]B�t�p������6n:V�_���9 $�@�p�KN��Qł�&���G����� �<����&<#�v�K7P��
ۮ�(W�����s�f:.�6���2�Q�aq{���+�($�U��,!ZQ��dS����<o�eNU�7���U�u�|�_��I����m�|�js�4d�tO����n9=',=!Bؕ��{.�z����}4�T��v��[I�g��e�Z�[��/��"!�=����L4�L�0��d]�����&�K�./f����ƶiO�w��������V��v����A��3��>y
9H��R�\���|�i\�T�C�:�A��k�ۧR�R�`��>7/A��Wg�1��r�8[V�� �l�~KB��sѻt����h��e%vd���V�	@UAn~wq�d�,l��xb����D��#"��$��PD���c�[M�ݒ��E���+�V/	�Ne��08!)pԔ6����>٨��օ����P��W�Z�!��j�K25�؈֛���@��+	�P��{��lē�
����*-���f����
ճ��rv)=X�Q�`Q�1#~Gx��q���>įW�jQ\\��-CI52���6Z�&��А�g�Bo��E�J���^�?�<�[��6�6�nc8�q�c�a]\7R�W�9ҪJ�ƎU<�ɡ)"ŷ�=��¿}UB���^œE�4e3�����.z�<�'HX�j��N�97 it���b�X6ׅ�Yf�x��4���%!�*r�'0�8|&@��;����O�Ȇ�B�C"F�@��e>כ����:�w�斮�w־jiW����W,�5�W�r/��Q��ǧ�O���Ҕ����U�7V�1&`��|\,�*��lI�jEt%ᑼa��l��py��نh?��@�-S/��y��8������LQ����󄢩3q������@m��
(U��r `��[�u*��$� _)���d
4�Wµ$����::�}�WTH����/R"'e֘���}v�Ziݷ��폄R�f]�N����JZ��V���ߗ����LʐHO��m{���
�Q��1"��CRR~O��w��i���W���V��QaRh9^H��EY<��IYB�F�(j��S�t�r_��D�N#T���t"��}���eT"��1*�YJ���w�~�_s3�ֱh���N:���C��YIm�y]�4�Z囲䛆	��-�Lr�L��:ɢ��J�㉷��b�^@���V����}�<�DD�4���_�
<��w�����UU����B�>_�����y�� _7З���p���CAi�	(�{n?��z�{d���v3�@�	�h;��ԄN�".�`���j3��&�p�S�[�'��Qٴ�@������sG��qf|Z��~�NT�^ws�ý�#�G8�Y�)j5�^(A���
�3���8jT����c͊������[	;ْi���ݪ)@6La�6��	�Z8��w�t#̈��Zu��	|vh'Њ�d_b�&A_in�r�&_��nm�U�:�����1��#5pN�_ͭ�Mr9U΅�5g�Y�Qq��ru��X��E��d���'a�h��ɇdO����)3.$>�>�yNA�����j�}G�f{��В5�]E�����h)��Ƚ��DC�x�<Jq�Lb���Ńs��s;�6�'��>PTn�	]�s�	��yy[���y�79��"��$��0V�އ�.��{Y�����\��wk�*E�Tr'��ͬzYX�����L�P�9�X
'x�±l�c��}yjH5���>Y�"|�8�ӎ��7R\V)��y��ռ�8����� "x�2lWݞ!���::C}.��t��N�"U��+�jݰbeL��L�LS���|��W.��b�L�}l���C�dė�ߩ! ��r�g�Z�AN�E�
�ϻ~Ub'|���۰�PJ��"R`��n��c�M�m�苮P���ub�c���� A�x�^����dY?`q"���Ӭc���z��G�`)�u��'�`���@X��}U�4���!W��@��h�ý�Q�N�Z���y�g逨�kk��J�xi�i��o0�jjq�^�B�y��" Lܢ;яF�ͅ���Vl`̷���������(+L̧,�ODx�N�.��	�"=N-��.�_� ͗&�J7�� �T�W�"�j�*�2��,�i��UE��4Wk�������2o��ۼE�1dNm(����9�;kGo�T�667$}�X�,j(���D���h��!��Lo�4[�Oz�W���T����&�1�M�k�k���B�f�`.Q�UÑ�',�6�#��-E^��{�o�2����ar����3��=�Z{_ٷ����
�{#�xk���{ 燂^��,���]T���T��51@����#�����(��w]u�4��HK] ����c�����ܺ2׊*r��9��.M�R`���nȏ���ax۲5\�}ʱ���)��	�n��{lj�`���oJWwX�;)���@i�'��&�+֏
�JV�~>���N�E�h �9d��x�Ԙ��I�%��-����%N��_�Zb�
yF�b���{���M�Ĳ�܌K�n(C�5�Y�lXx� i>�k�D�k�v��.�t��Q�@��i��b����-�k(}���t�h�Kf�W^�u��Fw����X�YH}@Pf�	�z>�g����k���>���qa��U���Ȟ���9�a�	.h��WoX��_���l�u��
��fv�6�RO��\L�Ho����M�%;'-=���F>�pV����Z-C?Z�{2{�ZE�C�t��E�(Ãd�z��GXOG4�ހ���?|��N��C�A:�90[�e�st��К= �\�;-X�5y�4����O%��yJ�zCC�Z���P���O�K�a��Ρ�2�6��y|~�WE��:�v#��;}C*w�$2"�J�􃢄'�(x��W���@��a"�+�R�MgҞ�:(.�f��jCZ��7�X�!6�Hˏ7:�dv��"A���4y���O6�Y´��g֜g+����ll��_���N��V���`��IR�ܧcT����i��EI�V�d���][\����qt�t>�%���l���N;�J�0�ꯂd͘�	����&��T;1�������=�}H�xN����<Q8����^Ljs0y{��v����t��`(��6�BKZ%��/b}p(�D��
"0F����h����]�]�hvI��z��[Q������H2p�yC����/�F�H �|�� �A�`b|����Gå�0R�b��m�}$]<����il�IlR��7%.�:�֘�þ�q�/A*��3�"��Y���k��솾���v���:����7�@���sB����+¼�W��\��	�~�
6�>�Fl�/cR�km��7.��-_��;��N9��0r��vO|��ր�n��
�<}���=1��c�~i��J���𩊆�B�/Rl�D=��ٝ'9Z��b��T�J)���q�d���럤��Z쫭8��r��%��	�,�ř�J�4�K7e��<��{ӂj�4��G��Y����Ժ]�"'2�ѶS���HE �́�ʯ798�I�&<=�M
�1@2-�%��l4�66&�U����T���m���#�?ںR��!(^�p�5=�mM�]�g������ @�������L>'1q>�Ī���O�i�
��㏶Q<���9��/�Y`xPQTT�\W�30,�X� ��<Dy���	�J�׍.���[H��g~ ؎�"�ҋ���0�Xij@#s)���={��	���A�tG)󒭋��>S�^�q��L��nBhr}0R�p.��=�,��$��ςd�GF =�:��5F����S|�x��F%o����B.�)���3��=�<z:�sj7�B�j{~�G\�*#ʢx@X�<�q������KO*{��� ��V���ƕ�pRϨ�������4h@�rm,��os�j����Jf���o��U�7"���j�<����;�P���K.��2�[�u}�lT��3#���#��˩�PNC���3\�@nn'P�����7�튙ܺ�:;
�����;��^/�o���1��ą��,==r�aB&�B�yF�3e6���=�}���J��J�,,+��{�_�V��&<k��+Ԇu�c���� '�=6��q��&UE2��Ҥ���C��xO���:�G
р�ϗ��~�0��cޗΟ\j��Qi���
�"M����p�L&��Ρ���	ʵ���s�J����������Q�ƥ/B���F`�21����^W>�-�F"��1�E� ~?�LB)�Vh�����^J���wsQq�Ð�r��!�֗�j��t:&`L��-���ȃ"S)&��쀡B�_���*�`�⨝����2&6}6�K/�����W�����o���g�7�$��ׅ�p� ��=A��ѱ���l�ڋ����x3Аq��0���7�)�׾��B%��u�jI�L":Z�5���/`^�W�Q����f�DX��Kأ�x7�M]:�11���M�K�6���Y|�Yd'�Z�@��`E4ھ��6�Ol�O�:���SP�3�'pV���*]�j8P���d�$�
��*�Q��.Y��j9<����O%`�\ep5'=��GX��a5�����y�2@+��o���˂��X����h�v��Ya��,�@q��@�b�9hF���+�g?A���+���\�ա�շM��"m�~ɟ~���v> ��$���$8���"�dws|���!���x����8��"��ߪvzꥑ����gR:ʵ��O��kcd�-�)U���j;	b'5+d'o��f����C�� �g�|��ڨ]=̓����:8��׍ Jg�A��k�o�ihy@�_��}��Y���H�}�J���:�e����S��%Ի�:+�ʜ7u�?�Ac�RcV�����n#��H�<�X��j����ᾖ
�ybW^��r9�M���C�aƨ���̗��k�{~Bd]C\���SUog)�	V�rl�A~�@�K����������Q���9~t2��^���.�[<�o�S8�%��c���]�o>X��4��8� vL����P�<�D� ��_�Y��7��[ t|ʴ�Vɐ����l�U(�����Z��I�,d�6hU��Hݹ�w�I�~���-m�E+�-�-�������� ��e�<��J�E�)��Βj��]��%��m V���~?=lUX�%����t�7o��G��-���
@]P~��)�4@���)+�g֟�W���-��X����@	P���Hc�6k���L �ڟ�XlC��/�.��-�6���m����	N����UJ�_l"�Ȥ؁����C*�b��J0Cl4��GzwJC.���B�� ��-������fm�1~�Q�S�3X�&�F4�S��$�9lm	�9��u�3<��U�ۨ7��g��}A./7��h�t^����s�״�@d���u�z�&���꾼wq�?!��2�]��1���-�>Ś�O�D*���H�ǂ=sd��>�^T��m��r�����s>!\^ww����(t؋E�p}z������tS��_Jrr�MN쟟X	��Ժ�3h'jI6�ѯ�x ����8��Aχ��W{m����3i*ݫK�IO,-O�#�3��{r쯠	9nI?՞f#޷��~���ɘ�d�vAl�d஖�7T���l���汼����uM8q�\h�JZ��?��r�6��^b�	azE!ۼ�'�p���0�Dojt��T�U_�Mђ����X-��%�����iR�\�ņHT�i��(�oF<��B[��Z��n=�Ne��F�!�Č(�+���VM�qF+Ar>B"��i�m��đ��ǩ�@1\�"hG���!;X��B!R�YU�<@:9	�/7IS;a�/}8_�tU)��Ks �8�����ZAè͜O]>�w����ߊ�B5U�>Pu�g�s	rׁ2��z8�����}S��sTˬi�dq�߃�ak?|`��P�����.#��
�^��b-�PGǶ��V�)����W�j�B-�[�噖)��J�� ���w:��|��C��3�ؐ=0���Q�`�6V���S�]DV"�"���tQ�z�aޚl����W�щ-��۴�-,�][_-�ԙ��@�"���y6s��b��=����>!%���?t;;���_E��L��5�5BN�#�7I~<-�L�/�[Ǘ-q��ɗE�OWV�
��M�dYLo���H��*�e)ÏT������+cP+5po�h�M#īӻ6[�q
�?��ΫPEe��i�c�B�bL��Q�>59��~62f)�����!|�PvaC?ռ�Ϙ�2YyH�BM����> ^��AD,�؋7���!Ƞ3��G1!r�<��{�6�|J�E�A��=9���%Q���K>�_�q�P��5D���q�����/�8�AB���Fn���ڶ��N�gg鈡�b�.V�𮌎 �Q�5�N��� x�U_�+��L�f�[������|6�+��G��	V��Xg5Л�ksN�F�C��l �p�1�Pc�h�$��2�e�U��O�GQ�/K����.s��gO��v� �$�O�03#��,Q&͚�f�]_�B|�����~���u��n��V|�.t#V����n��V<I���Ҭ)�����7I{�RlGٹ�A�e@03q�Q��Bb(��p�XL�jP/Ս��̶��Q�Bߔ��W�K�K������g��D�sʕ2��$>CJiv�aǄ��݋�Y�o!�\��ZSn��q �iPZ�;��\�=̺к���/<�|o8�v�ͺӡF�.F���i4�L	m/$��Sa$WK�ՈP��<'O��H�<JU�C�eg�:���uq/"��Z%ݘ)�M�C܊�:!<��V��@�ت
�s��E�Q�u1���.~�R�����x�a���������=10`��<Z~ۻΒ�}��h��ߘ?Gh)����
+*�g�Z��)��@��_
p6�>�4�?�?�����َ)�`��gfɵQ�c6���A�+H�����t9d���R����b���Kє�c��@"H�>PA��g�ݟl9�į�������x��Kx�!M�k߬T�1��gk��y�`9'��z`Pź��A�����&_ ,�a���U����ڰ����*�=U��C�)�j����^a����7o$�ֽ�V��(���ic J�y�4�7fz5��P���G%��^S"5 �W 2���w�� B��ݶ�"ө�㳰��(��Fy��Ɂ�[^H�S��>���M�J��|=H�!�:�i^R����X.)�&�`;�r���N6�����w���×�*p�՘0!��F+c�c��yh��.�!�EN����Y�hc����@�ͼ�
�h.i+5��H^�y�PKJ`򮢓5.O�r���B$�:@�[d���p��t}�B�4S�F+KX�L�96�� ̯�v��܄�o�h�����c̰�y����#x���d�����d?����|U�)�r���r��F3x���חQD�Pb��/�k�eِ���p�{��;�s����S=���Y��(Ak�pG)�_҉��%q�'�V�O�F�
Ad�@��;�3R��>�{�V��o�3)KT��H���(
h*$.|��
�<ގ��}���2��~b�#-E!�Q�H��tq�L��M�0�XM��֊n����O��v	���y	T����+Bڮ�?�"��aY"s��w?�t��.�.�Y7Uz��d�����a�_"��.ό䧴�w��=��ޠ�@��$� �j�
�̌�w��3�}���_��s��H�W㥈V3ǖ"���(�&1�!pB��Q�<�hj�4������2#w�����ߣ��yu�(�'k>)d�]W����2��2��UϋU������]�4z?���L�� ��Э���Q(�{���A�Q�ܜJs
O�	\�KLC�\D~�IX�� Wt��7K��(�g���y�'�92)S�d;��g-��k)�s����!td��*K/Z�Q�,
��jϧ�$�b�a��������������z�
��q����yIx��j��@ܙ�w�2������mQ�ְ��K?�8��~���ΏGtK����b�-�Mj� �7.� N���G�Q�*���7�魍ݾ�>����ȁ��'�����n������~�����n�%�}�lyS_H����$�p�wmúu��X{��cZ�Sj�u���L����{��5��#c$���ጷn�ws�i��'j��~|�h�S����3�l'��hG�����n���4G�#�ec�H��DM���C7¦�[�CV��8Є����A�B�~����� U��g}��2��v��F���n0P�Ϳ��8����3��=��)7�>Y��ȫNk��ܕ�T\����;�4]���ݾ`ի�j���X�
�R3X���]wpsb���N�D�Mm%�z�a����*V$�ԟ�?�bL�RRa�}+��a�wB�_�Nݧф��R����=����� ��e�UR�A+���8�ώ�UӁ���Z�P��h�q�,���
ѵ��z�iD�T���ɸS843Fn�P����N�9����S3tx���x:� e�Gy����j�?m��`|���o����d?��ֹ��}��a��t�zfBy`]̋���UNd> I	 w����/k������� �iGI���i�Ȣ^UyهM� [�V���ˆ���������]��ʼ�8�U�U&�#��!�
�� �K��S���eB̏��������]W=Md'r�}��?�BT����Wv�3�9ln!)��D�X�oж>8V�e��� U�<cA'[�Nj�S�:��PXc�]�ϸ+y�1���mv���CQ݈v�%�sn��M٧AV��M6�3;c 	QΑ#��t�)��p���Fx��j]>��8q�C�HR,6�q���^!�0e@��i�s�f����@�<������q���PU���y?�x��G�\�����G(|̄����.j�7���e��aT5�h��Q��wA{\J�̋SB�D��2 ��l�t	{Q�yO�sj��3L�(��၁S�)S%���=?:�O1�Ж&KǍ��my����]��"�#6hĝ$v��a�΂9
����
�Mx��Vj�����y>���^E�5L�����q���c���~��;�]���affx5g��'Y�����
EY�����&^�ܥP͘�X)��f9�*����t"�UK�EM
�w�揮�5{zH�S+3S��R����Ie�]��J4E%$���G:���7�@c�F�I���$\�Ã���v��&���b�r�|&CA�i]R�f���ѐdœ�0nm�����?���BkIXy䬫���$d��Ϲ�3E�꾀D7k@ӌ\f6I��~�����c^I�d)L���u{�w���N:8��*jD�,��Hl�?I�d���flv��l1�e��_�O���ř� F��*�D��\<}O�b�n��k�`J��'5�|��LѪ��l�T0��6��y~��<�W�N�Wc�W+(�d�*��g����+83ogA���2�3[�;b+��CL/����m�St�&6�<���̦�x��3�0����4�UGV?gU�/�{L��&v�U�Н�7��;�?��)69���e�����Po���D�@���%@j�݁�j\�0{����׬2�KX"�U\��!GJ�(F&-��|
;& ��e`����t�׍��of��+c7ȃ���	k��l���%Wظ�	�!@noŪ%]��Sڊފ������%wo�N������;�c�����j���!�뽣��Fo������}�xUK�-!�L,T�>Tő	���ՎO����r6���-�F Sf���6���9�]�3Y�^Ut���m��ۂ�l��0����ꎬXM�1�&�C�/}	*O��ύ�532�qd<��hT.+�7bR,����w�� ��3���=�����H�(� x7"$sh�Yʷg�~�ъ���ǻ���9.�����!|����3�2d��O>���［IvG43�0��U���L�`���� �q/�Ң�b�����t�a'�>B�>,����zCn8��aƯ$R���z^P&y�Sc�ָj��c[l�'�V�^Pk�o����ʠn�`�^y����Yds���N�Y,��	D�;F��`J]x��R�ϓ�W"����a�%��?���C	���{���< GƘ^2.�T ��nW���y��f~P�e��^-v��-�i��"�CT��4�mRR��rʚ��m�&Zo�mڋ��1��h?���̡���D���k+*��˥`��(7q�m�X����+�m��2Q���e7;�� �n�h�#}n "c> �-]Z���>��5d������%J�`S|h9�b��}X.+E`�h�ɳg���2g��$�|�<����k�~R������8������� �Px�hZy>�Ľ-��j�o�(]�H'Q���&\;������Dń:+�}��Ŝ�Sz�|2bR���l�U}�9	�;P_V��4f;�_b�3yXP��^T��!e�R)a�
�i�؈N9̓UM��d�� �;]��-m$R>@���(82�؛P�QE*co���¶"Z����O���C��[�q��7�kو)�M�쿘���w��]U�ﱯ��6��^��
�m�f�+���E��^ń���������e��$�/�{M�����8ig����Z�w�CN�Hnp��F���Ɓ&4��Ұ^��$C��	T���3��K���G;7l7o�{�#n�|Jv��s
0��7:���Y�8CVfke2�\.�E�wᳺW�U'V�< ��L��6nd3?$Ҳ���pq<������Y���Yw��T��]TP]8��^Ev��˩L~��������.͓�v��������l��[��"w+� �E�Y͌�W����j���̧��M&�<ϔ�6�߱23� �C�����LG>=��r�$41Ӹ��{�ng�W�ܧ^9�����@ҭ�h���v*���Ɖ>�7W��a*��!b��@܋� �H�n��K9_������E�s�@3��է=��fy� ��fE�D�+�a�e���������K�E6�%�y��(��,O>e�Mk��W]��~ش��8q�ݍͿ������<����6�WN	rrh��Yg�n��1�.&|��噾�9)���"���-cq\�|.����7	N��ne�y[�ڈ�䫎��⨋����D������T�Y�B��*�޲4E��oz�L�1�-�}j�z���/�k�Rb{��� dh}�M�r�I��� �Y�q>�� ���?�IP.ትʕF��nޅ$ÿ;f�ナ=�*��;���c����2ˠ�����*:P�Ƽ0���&]G��8��c����Ex��F�>%���ʫ[��Bq�%�f:������}w�'��ӎ;��3!��ej�-�2�_5��(
}�oj�	�3��v�a�V�!W�Lu�!���4�5n}_W!�}�!d��7�^j�a�Y�h~	��x�A��Z��E�~;�D�\J��\��H�����x,�w���7(~�F�!�ƕnG�I�ϘHi��X(}���>Q��z�����6c���F�:�^��O�)s
��]xHcӘ�+`E���yJ�(�L����\�s�?�6�5��怶�����Qψ
g"��F0~�`ϔ���Kk'��z�c�|���?1<�I�����X�g)]Q�C��W��g�A�K����aUW�9�U���sv�� ��OK���X� �Jc�_l5k�7�n�b�{�?�X�;���C�^S��To�h��a��ʔ�˰��~QZ;#�~kȾ�1��Zepd�x���y��u��C������{��Ew�_���lu�v6:̞��Ұ<��ղ�7v�:&{�µN3��Zs��~�Э�H��C����i� �AbټWTl����G��U�'���(v�)�惮hš��N'?qc{�h<y=ѓ�eN�-�5KyzkʋIL+��u�C|l���D\��g���jTvS����b�	')r������"�  ����t�\��q#��KB'�a1gW�����w��{ {�I���L�C�B��v>5���y��N�1� ���v�R+1����:T߼�M��1���pt����2��udP����(8����DY�e��>��41�o�n̚�;�l��?��r��ʫb)�[�g" ݻ~1�:9b�7�J=k�������u�>��f可������"�$Iª��~T;�j2�&�e����Z����m�;r���f�]��f�5s��=|�D7�1|c�@~���å���L5�i3t����f���(�)�0��j�I�ޒ5C5 �\�����@Q˯4�^)V�����:��i�m���`Y�ؔB9+�QGKJ)&1w���ߧE�����o�k�Tݤ��,czuq�\&�u��B~'���jY�����5��P�'߶�����QiM��M('P�H7"<��T�|٧�@�����	���ٹ��h%v�Ԟ	�4�8��ːQ|
����6?%�	�M���[��6��p|S`�v�\���z�2ƣ�~L���/��Yʜl��L����m�����*�/�򀚳z��и);�y OU���q��4���+]�ԽʼİE���9�P�`� �s�O�T>�H'F)q��.R�����ј���r*fK�AK@�R\-.�	ۡ*v�R�o��a7��݈)x0z�����2Յ�\�l�x��f	O��ң�-���=��T?�ͫM4�F��lJ�� v�@���WƆ;є�%�u����Qz`X#Ⱈ�R��"�v��E�"����*�����ڿ
Ql���^H�r� �F?�'�=�i�8���h9�d�Ԧ{Y�!t�uת���1%��TN�������9�&:+I��M�3P�����$��c4C�E2g�I
�b�`O"0�J`�'�0 g(���5jލ�� � ��k���C�@/vT��Cw�R� ߟ�0O����K�3���ؾ06��^{$�a�q���7s�n�p�� ��)(�Y��;v5GP65"iB��(��~߁�˿� #y��X�/�-�q�����$���������S�k�pjiȵ��i��JDFw�!�P��/�a2BMgHG}�Z��JTa��6��-�_�T�h=��S�@�H�J��pS��Eu��V:�-�
t�|��O8�8�#�G�u�a"%I�qwee`��Q����BI�@M��*˵0¥� 7���j��[#��I|�J��e��'����:��9/8�{�q��6m@�7TZ����B�C�������m�~b�Ԝ�5�m��`s�p{.���J
o����U��g�0An\7�#"s|����t.�WR�D�7��㐠�ն�/C<[�]u��(��̾���5�v>� ki# � �4�f�h�����_"��AX�4E�\2�N�����1x(}"C��������4�� y%�V��'^��B�Om(6��\ab���'U��B��K�\��������u���|�u�n�!����XGb8��[�49/T���TaqP�G�7�*��9F����EW�W��	�5:��ƶ�[�|�|߫/e`SJ/�m?N� y�H2A-Fڞ�><^�בMz�B2�3�_���e��>-�x>r�-yg`���:tT���,\�u�mQ��?�=htO�<m"�:�Jup���JV�.��5T^�
��󄦕��x��BR�� m>=+bڭbK)@�Z)���R�+���'�,��+T�8��EK��XB�<����D���b�!���$9�O��k�>_�̇S�C]z��A�'��̺K�q�~*�s�`�k0A�
]���x�^p���p����t�ps����8Ȧ�T*��眅I\�?�[�Uw��T�~�O`�Ɯ�S��~���������V�L)����6>�\�
��h��w�X��7�f�ڠu�u����ҹt�ɥ�r���
�P���nx�
���n�x���ܢ��u�Ћ�n�7�-�[]K0��!b.���l��ֲ���eM����"}�U�Ɲ3����-x$"n�<{�>O\UV`g���]��b��;2c�L	T�׶��[�RYM� #ุ8X�`�],%�ׇi�T�9��#ق'p@�AQ��W1޲��
d  3�
��X��HAL�Gb)�E�|�E~��f�S��̕0�J��S��^,x}��.����{�V�?\,��Ǹ����C!����у:�H��4K��P|O���lj�)tY�����2
��1���"�� 1�\���L�6��z��{���9�42K� pX@C���&H72��\�0��$�U�e}K�v�刯hE�1Pdk�wḯ�Ҝ%���a��upfĵ7̤Z�~��o��:���w�;q�0���q ���:u�#����m�
ʟ�}��Ə#�<CPT�(X%��0�:�ē�E��ջW���`��$��&�����w�����z������]�}��g�鹂�Ʈ�LO�A/+�(�+��K�3#E�����Y��sU���L�=�P��bf�z\g�%��rw�dq6t?/]���E�0ڿbB�,NIa�w8�Ԅ���/����]�p�V~�gMs��B�F�Ӳs[�&�ee�U.M7��"t����q�P�����d$;��#�0��I��攱�!�֪�e�*	�o3��~�:V1�JJ�
���vn�=£k�f-GjHJ�l���u͇�QM�����\^`<�7�$)Z�(0"�/7���
>|���4cJg�.l�&�&��H�;mk�)(�%HV��zO��]=�ב�\I�����<'3�Y=β���{j~�R]gın�=
��P����)S�s�eu���'�8�\�y����zI��2��|/�'���%�;��,�* y�.g~�+��i?�s��\Q�]�O�����T�<R<��K����=!��,!�a���<�0�K"�f���9�A>Oa�pw���Bq�Eå��J�#�3�#�D3��9k�.:���C�z����]�������rc��o�G�;��0��;JuQ,H���MA�ŀ�݀����w^�w��i\���I�q��1
80>-�,M�Vj��
UK����@�$�癰��1)CH�0���x�\1�4d�`(~P�03@yOˢ��x�w�"�-z�r�G.�|�g�D_زkM�|��'0�`�'��Qx�T�K(��,�E1�<v�H~�<���c�ԑ��Lr�C|,� �6�K�������A��bh�,]�8�˴��,���l�B\����]�؀"gz����
��X�Z_�
�o��QM�c�D���(��@����1p:����4t�A����؃�8��t�険�����[E�n`� k�O� �k <�Ή�
H]��z��n�ts�,}\��@1v!د����;H��?��d`�c��b���nݨ0��u�!�O.)^YƖ.ya
E�[d}z�j;ÏlLюn��ʬ90U��0n\��S�ͯm��P[�ֵ?ݴ��صs��6�ֳ��J�9s�N�����A��DZ�����g���cA���N V��۹���;����C��*��������CjE&θ�Q�r�X��f�l�vI8$�6�<��CZ6����:�I��0(��NW/|��
��(�w[D��">��E�31�HΣ<nF.��B��i��8X�(��[fe�В��H��T:� i��ֶ�w�!P@����?kv�_.��)��&�:�����@l�i`���j�R�v�݈�����=VDs���w�$\x�(S�*,���k�.YrD���E��Jݏ��ēང�:ߵ�-�@qT�}k�KtՃ5�ZX�%8�R��X�u
�s�}�^"��}K�K.����v��	�4�߮��^��xX���2F$"7u~����F��V�֩r��{�m�g��G���QL\��6�)�0�k�5F(��˪��Q�Z$4�{�ɓN\����{�%� P
sY0����w���U����uB3"&%�IFR�J%�8]�D�ڻ��`�8���ޓ��-'��HUd�i��\ͨ;Dl��������g��B�#���*'V��S.���4>q6�n߹�U���3�I�5�w�ё�Z ��I����Ƿ(�(�z������I}cO)�P�@W�a�!ռ�OQ$�Ubm㫵S�[\UܙyuW���u!�C�Y%���]�Z��05$dq0e�(ϐ��0�j�;�l���/�W\���dУ6�ʱ]��U�a�l-&�I���-�ػ��h�Q�Vc�,����j�<���F=7|�ʙC�
��7�D��ǳ�C�� �'v�m�-��P�W1ϳ��ՙF�;bD0=n��
�AHO|��w��0����@S�d���V刳aO�x��l��Vծf>�61�E%H~��Iv�JF	�şO�(�$䵏�rz�{�c-kُ;���U�y�"\���4&�3����M�eH?���7��z�'HI�f�s��x`j���`* h�f�j�Z<lx��P%ATv���쓲5���7��F_���f���Q3)��~P��Oɥ%"{R�Q��|�O����\���Kӧ�'qv���i���d�$�;�f���ː�U���w�w��P���O�,��p,6O���M��Z��/Ȅ������g�}Auk�XN�x�͕zQ]+bO|0<��G���� r/��2yQ���.q����7�Y3�W��uk���~��ґ�i��z���Ճ� }�����\�`�sg�[6O��ެe'������mH�l�����$/��e8ABx*L�������0�9eϵ!��KfZ��{�D����{-�{)��`����?���a��~/�W�rC�Oc�lo�̉%;����^�~��%�-�b6s!?�3h�\xMJ�,��ҏt��S4�xC�K��/� �B��n�jA�;��w��Q��R�&4����/K�"b�.i�"��9 ��ǄXmt���Auz���v�ap
�3��Zd0җ����z��3za Ň �L[PIs!c_�h��f����'�����8����w�" ���$�B����6�	Z(r�$&�Vq�;��ﲊL��Rr(�GޏgJvx�C=B�;^��m�m��̜Z��U�R{�ISަ�΅�v�4ĀY�!�4G�*Y�އ��.k1��������l�ob#(
"K�j�40g�:�)������C�G��f<}<m�	_&��8���R?Y-�H�C������^Uޜ�"�A9U!����CT~��~iڕ-��k-(�'����?�$��jW�
Ρ>W4Gbہ�0�����Oe�$�
�bou|˔�8��p'kx��=8Qm�K'g�S�ZC ?`�x�Z��8�����	Wb�y3f%�DN��Җݛq��t�?L�O�uk0�d��gs�Hb�tH�߿�Z��j�o�����t��̠F�������G��b�=���J���*A�H�m�����ƽ�s�(�mmoO�x9 ޼SvU.���!�S�A�P6��	��b�6Na���"��YSF:�4PRէiq�,.��{.��ep�����z	}�fK����U�r5��F�2f�u��*�b����G��͊�(���Q��EE�}i沼��xF��"$�Dz<#�XS�B���Y��8 .�	XQ�SV��Fi^
2[$_�ʹ�0�##4��~^��!ўS��jJ<����L�;!7R1P+���ĩl*9�� ��F�Hq�
��$
�Z�?seH]ؙ5����~����}w�kUg[C��_S��s�N��B��AQ��	s)��1�^�j�JK��f��O�F:�W��B�
(L^֥C�<y�`����QF�R��R�������wIe-����:�H���s�!&�*�5��N�ɯ�j�Y��z%�9Z�r��Q-ϼ?WEa@��X�ك[���~)\ɕ�gX�|��.JD�j��9^0Ծ�ZC�����iU�DY՗��2�K����W\���oKF#-����kB�`qfZ�ښ;���i��3��fl�͋��J��9�{P['���j����P�N��)�.5ԇ�����`=g
l���V�I(��u��0(�s�Vƍ0�`���k��Qq/��1���f�FIڣH��>ʒ�ف;�i�a��r1���9�QlS;|LR�5U�k��Iw����}+׾��6R^��ls�=�2K:[��!��wR�{pjr<�0��udOed�#V򶇪��W���y@۵*�����}~��0����M��<�Y���o�Z~C�C����/�*)�5l,�.;&��D���e.�t����g0�#F ��G�$�Bp�:$�J���h�������6��tILK�,(u_�֔�j�U��7u����>^+6�"��v�j�.3�4ͅ��fb&Z�m%Oh�K�=���AE�4��Ᏸ�K�p��,1�p�Q���4�&��@�U���c��@a���<�>%V�@��?�&�-P��\��- �S��b�� ��� �S��x����|��C�ӎ���I��=����H�, t�F��o�����ߜ�.1�"d�[�<�Х���6��1�WD1��gu0�
x�'�;N/r���'$����=��i}�`\w���$ �R��3'W��ؚ�8}'ǆ)�:{��@	����(������p��-���b9@d]%���u�[{�B|w���'���~��4>����j�6�^��T9z
���Yn�ix W^���͝�.�b�T�y�~��SF-�ia+!\��g!�;-��؇4߀�s��/
����Hy�=1����-Y� ���$U���.\�|���w�7��q�Pd)^_,S�@B	��Ӌ���Ī��'�w	�m�N�W���B3z�ׯ��:��������U��ji��� ��w2�P��}ٺ�e�^Z��)�s��������>a��q���u�V��qΏs��0N��g��%��G��7d�w�3k����0	��`)��k�y��y{1��}��M��_����u�;}H���=U7(�lVۈ������P�m�3n:����Q�����F_t*x7��<�F�mzu� ����Y�^�տ���3%8�������O����b�ѱk�ؤhxB�C���s9�~Z�3A�ƀ��8"qG����)WϞ����Ɗn�sZO�j�G	��f�1�Pdc�CT>�Q���'s�\P1>����^���l�{%Ѣ"��|�lɖN��G���e^�x(�O��1��}M�󭳷T��oZޣ��'?�o��9�d��D�_&��)������5�ţL$%�3+�5P
h���RI?&���N�h��3ӝ'@����b�|��D�݋b��NS�t��2��X��Hsx}�q!ˈ�W�o=0Hј���T�
'��/��jb���:�������������.q�1��ݥ8����`Y����,\�-N:G���5�
qO	 � qA����F��_���e����1~�3��2a_��''X�w_w�R4B�?cn,���E 'J�8��]L%�@ebe@^�G�Wu6*!7`���L���f�(��l쐜�B��B"��72�$��b <ʲ%��l�Ʊ[�zʦW�ưD�?�F��
�����,� r���8vU��0M��H�L%*�7Z;)�Q�}(�V &�כ��?�"\��dÇ�&�؞FP��?�A�ޚf>_�d���N��m�w�Ц�YD�j�6"%�{�N~���~���!�]"��Qd�4�H�;�$x����Z�r�aC[{$����/_q����v���'�Sz��ͅکq�`-λ�͇1��6|*� s�,�Ύb����ٔ$�qǌ@�0��={��-z��կ֨��k�Ҥ��u�YL�ا�Oz�����	G�OٚB��t�O�"��޷��k���"S!y�i�8X�7g%���_�5.�R�z��"�p�1�;�`'g3f�s��	�0��.�������'i���-��F��������l����`���?C����5P�Nː�k�+�h�>H�ɪ�V�]��u�j2�	aXv����t5�TZ�+E�D����KԔ�a�� AH����x��XS&/��>.nH��|k'�=�3 d���?G�>�TxE0nnJ�v�
r�v\w���I���r�G�h�br�+���=ݪ13y���e�P���ݵ�IM�v�La,���p{���y�S1��'S 2s����tV��?�����8���X���G�.f0��P�GT�����'V�ꕚw˲ax`���m��`��Cz)K^�+�u��b�i�m�p��#MM%�Y�A��F?�jY��q~���$e�D�,�	>KE��7r�i�
'>��:�R$J��JH�W�t�:���W<<���]��"gw�Na\��RO�#n�8M1�Δ��F��֡.�N���F%΍v8
.
�"{�p霢r���Qĩ�0ʞ/���x�Wh�A_$$~=���Y��P��r�2��6���)i�>hh��4)Ps&9 vW���c��l�]���;�_K(��'s��I-��$�yjWs��SP���f�Ա�py�[��F#��apc���E�W�N�rG�N>��BtS}`Z�n��]�YbEqvl��L�Ll,�_qO�H�PZaަ���hҽ.^oeĳ�Gzq��VM���5�g�<ڻ	�>ڑĩ�dW6��4�1߱`Eא��f��2�(�1�-c���ύ��n:'=�? ��>v(��y�z/AR}�Wc,�E�Śr��(#�EM��-߿_�d����r,�xF
wH6�ݗ��=�xtz}�Wer�����r.Vu����9a�3�n�����Htr��p�]��{
�;�"�RO7�֣�X��>�Q�����+g�YU�m#���9 �F�M�o�xɎ�aY:��a�w�'z�@�ߦ��C�+���'ב��z/�U��CSq�h�,M+��f)ˋ?!`�P.��&D��5HS9�p'X�X���9A�J�v���H�	�MD��-��e���h��x�d���J�Z��`��I���#�#1�����0J���d��AY���
s�%U
H]� ��e����8>RJH�u��S��d�3Ҥr\�$�4