��/  'd�N�d�}���ts6}�>{8�V>@�<a�4�<?���>\�.�"���׺��Ie�rΰ��g��j,�N��>AT�<�X�@qv m�2 D	�	�tAA翭�D����v޿=�\���.�"b���J����\�6�B36���4����sOQ'�B��nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n��:>7ߎ��Ғa��H�Ɯyї^sXz�1>l��^OɧF�e\p��.�Բ�O�mVZY�5FC�l�U�B!�ZZ.n#|��}���{息�}>���� �������U?�1c��Q�����wKp���m
Ǻ�F��[sV������ �J,a�"�Yel-8Lz�]7�;(�����:�aOj�'�0�X;RN��<r���M"1��8I;2@]��,*�>P��Ƃ�J���ڊ�;�&G�o|"�����U�GX;=��#��ϝĔΖ���k��U��A^4#�����=93>�ϰN=�_��}I�v"�{��ňR������e�k~Gڞ� j��[�oޛ��;82{�;#�{��@�iL��'�7��r3i�dY��� ��i�"�M�լ~[�:х�0k�!�g�`�n�L��q�<sm�K�kt_8R�_�p[/�5t�8C�ӫ�b�~�e� 9"&n�i&̇��Kqj�>��
U����ğаV�S]II�k�ą�?���lE���4�>�7E:��[v�:�pR�����U�qq�_�����".E5��@�@a��Fw�*��R���J����)��5n�6����8� f�Χ�E��y5��p!�����F��6�>`ä��h9��9ΰ��W��`�xy_��|��a?������a@�a�U��9��E<:QǶ��.�89����{г�^ �$����l���s���b�oI��}���ː��ഖw�A���ܪ�h*���w����|D=y�|�M/׶�zA5�[���?�Ct#�Vie=]�:���S���?la{X[0r�OX3��H`�FCq1�`�g���A�;3�&�V���R����d�`�.����zTWZ����B�&qǫE�~�jUҬ��&+����! �~�J�L�J�AMPs���^M�]�ڨ`?#(����J���y�]/Xj\�a�n�7��/��
�A�=�����2P%�
 B�L�V�Kl7c�S�+;������u=XJc���]��~��c�M%K&��V�������E��\�i*.
�J!"��K��L^��N�/�?2��iD�*�ך۹�� Ai����6\�s�����������rm7�� & {cr~�.�j��"��l��K�^׺8�_�)�ӝ<X��3͚<3�Y2;�$��]I���[M��)(�>�kb������Tpu�3�	ѩ�ʟ��f #��"���P�!��RkC�1Z~�_��&�^eq��w��W[X��I�b2*�q���ϰ�Bp���������K�빻p�T�>�b�<C�ۮ����^1�&g8~�$/+�����a	���bc[K�ym�1=7=ջI��|_�v�3���� ��̓5�nP��G[�%���2KsO��a Lw`�g K�����TŜ�W��0 jidꪸ<בX�^b<�*����4n�s�Q���|�,��z���U�c��|Y�oS�I`N����I���2t�R�M�����-��⻶��I��}<V��܇fB4�,��a��=~����u.-y�d�_is��J���t��ek���c�����ڪ�=��z���\���c�?*�z�-�1�;��7)��3;���{������+�|Z�#���QЙ�A�=�5����Z�\�@Zqt�z,G���4^�l�<����}���]1_NAyb� ���	vE�����cX��t�/�28�x�̀���v+D|Q��ňO�Lr���{*�Q��.�`�&m2"�mZU�G��F���h�dE�љ�*x�5�A�w�U��d%?��-0g���F��Oa-�7�f������<����u�9͉�Ľ����Xzu��[����	ufp�f	$2��k(�Sa�����J�?�mi���"
ֳ٦<{����A��d�ܳ��$Z��������S���E>#5��W���S	�MX��jð�Μ3���8�q:z�.��������߽;�Y?�v�@� @�L��φ�M�hV�r*��
iuW�@)}>1L�w��) ���O�%=��?��prW�YaU�����*��+:遭WL 9V�D!6�����<I�N�I��H:���Kf������a4p\B_�")!w	�(�%\AT�������4�s�.<��6))�4�2�i���2z��q�/�͆�}_ڛ� (��>�����Ȑ�T-s����j�>��^��oү̂C��lF܄+�_�Mcͺ����5�pE|�o=�(�|!�5��|��]�!qC��[v0S���a"H�	�����Ļ����!��(�]9ϩ��Q�o���ҵ�èM̭f�Awt��<vU�)N*�u-礃�-q����g�쩖,�>�%-+���;�l�PP�I�֊j���g۰�v�DQH̏�T�WD�A�k�A�^����7�Mi��� ���G�7�m�;ّ�f��3n�W_�.F.��t� ��;��C(���h��a��޾���hz�Sm���m��W���{VtO���N�C���u��'��F���yi@�qo:LJ�SЙ6K���!�t��0!
����4��9ztM��MF�K��P�� ����1&������bj��W��o���B+a$�q�X�7|�\f��qB��k%��ȱ�9��b�)|��%��1�}��ڦ��Dm0>�#	�i꼄r=|�����r:�[��{C� &I�����85�1�[p���`�]e �x�I��Ƈ���PQ^�� 6�W!J#|�ea`PEJgt<g[�	�+ �x-��ţx�x����f�I��9�D�ي�؂ϸ(+��	6n�#���?��>��Č��л,1W�|��}�N�W��R�$�w`�� ������=�p>�Re$�p�Q��p����e%���������Tg��;J%�"g�p��{��y��R:��U�*8��fpLѹ [h@���ms1eKDj�+#��x�9;A�}���d-�u
�2	��[�ӣ.��D5��:k��ld�{T�n��M��y�zd>i�9�����,���@�8-U}O+���+w��Q��jS@�~g�:GOW"�T�7��H!�&L�
���U�C���(>5!%��S�To#L�
3�/�Kfn��d>n\���$���\6����B����4uڵʤI�L�a.�`N+=��@�C���[���N�ơ�(pp�\���b�͔�M�cA�1����k�%fAԄێ�]������+H��3)��f�`�����C[2C�Bz�V"��(�|K�Ə������kH�{��r���Zk�"�%4�i���;'K8������� ,`�W#���m��ނSr>����7i���Dn�ީ���L�EwUSi�a~��'����EA9Gf��
��-ӄS)z�J@A�ɫko:I�zhZ��%���w�g�at
)�O+l|[�Կ3d���j>�94Ǜ>4QlM������_0�Z@+�~�+�|ۿ*�ԟID����p7�r���3�uQ_hne?t�Dp	-�\�#q�z���oeQ�s��fe긥���-C�v��vS��ƻ	Z)����m�3� 7b�9<(p�κ�=?l�~�B�.uK����%�U�M��K!�k���up�s<���;!���<�K����{A{�Y�ȢY�P�l,g�S����ck��i�������:r�V�Q�΋��\�m)�\%��\�d���["^d`M�o5Dp����&Dl:A�$̱W�ч/�G��If���V�$�Ē��G�˶��S�������-�Gxc5
�h򪮵f���ඣ�-�-̲�S]�箣M*Y]w�P�k�)��"�˻�)2l�+�7�Y�b�v(˺�u��S�&4�G��G0��=d�H��w#��
h���SB3,��4�F���GQ�XI���u؃�w�����Dm��b�8h&N��m��Pڞ�?ʟQ|I:��o����
�[�f9Q�5�DT`ŉ�Ǚ�'�>��l��&���%����}�J~ �%�	Ē�ht�8Q&0d1ӏ�w!q�w�>�I8��+���\�hs�]�sZHXU�}�>�`�T�Ņ�vxk�p\������s敤Jo+�M�M�Հ�>�J�<W�C��ﴕ�޵uf��l�u{p��-�^�ޱ\�dճ��[9	�v��k�o�H$8����bU6�l7���E=�,��}��w�ɂ������R�q/,c�bؚ"A7�A�]$��MqG!3���k2
#�R��B���VWQ=���Y��l|D(�'B<�fTW�������TX�/�&`���"6,CĠ^�V�p�$ۖp�\/���>TB�Y�1=�.�I�^����7�����T/ʧQS��Жýi�J�E��ޓj�ˀ��El=Ӫc��濰d��WQ2?F����+/�.*?����V"���|(�7�1���K�L��Y�O8��\f��z]E�C(`�&�"d6a@�J�߲Q&�9���C0�'/�z�ov��c��݃�ӷÝ����.�o��S͝���h�8���h���d�Pь]h6Zo������ˇ23vo�����/�XK&i�|}���u��c�HW��; �9C$�y泭���l��l&��G0?��_(�||%	x���X����k���E�Cϼ��^z�I��u,�#�@p�</���۩mm#�u�4eғOG��5��\�|�U��� (Wm^��Ev������L�5��d�,뤭M��.YN|��En�28Ē��i�7�9��R	a ���Yiݕf�ߝ�\�L6�����<?ss��>wR�Q��	�RBi��u��B��`��|�@B�[hX0 @��(���EC��x��qaF�TVr�a��ɪzHgt�Ƨ��`���).s}s�d��o����(��xr�С����X�#�q&j}/��n~�m�0�&:V�qz8+1�n�9;4����!��r��4�~:
�B����0����u.�;��fp9{�����@~Z�!^�hC+gZ"~���I��N�+����A$݀����c��N���tW���������C�ƹ�1���Y����������)"���g�䌮��:�!�n*K�S�l�t���]���cż"[�y�N�%���}��1��M�6ٱ3�UT�,�ה�A�6�:	a�瞾\�|[�Y#��;���;��z��w���ٔ&s�����MdL�xu���#	 ��}?ng���3�y�C;i���W�I�����͘CgTQ8+��k�`���[S������<���d��� @�G�7#Y��� � U�*�-yΆu�&������<Ww��ͻ��_�O��cFH�0�=���0�ԋ��7CE��HS�lC����	j��XɓiҶ���A�zVv�A��C��׵�kmT�;�'�r"�$���lD%��)��ׅd;b��.hJ�X����u8ê��ո4�"A5cߖ{�{|1c�O�D���3�k�&��3��pB&U�˸_o[�Ʌe��*&�kiz,�T"�2#.]��\�ޗ܍�*j�Q~� �堢.���p{@1GZǂ��=�s��V�H�O�f3�ok?9�)�;i͡��o}����n��"ӕd#؝�������nP��to�k2��}TE�H�D���د�@�.tQV2:���U�f#��[r�6����#��k����6I�+8�i�U[�&�v���u"����voG�����E�"x�����;_Kܨ�gA�|3(A��L���D��#�Q mǻ!������#���ç>��3.P����i�;$�q{	GN���*�^7!����i/"�f�6�9r���15̷TqK
R�$)����q^^�Ld�9��t'_v{�{i�f�#���`�p,Z�C�Ѱy�t�ͪ��$ �_$^���@<J��AZ���yqF�OW�d��PE��:e~4��hv����|CT��1�$���L'W���3�~�\LaZ(������ŝf{�wE��&|{�����]p�kb�Ϣ(���k���TϾ?w�$Y�1GK�R<��)��6�RjKOn+�|�Cdrz
W�Z.G0�Ο%7��C-�v���ߺ�<��#ziz�=�����w����q��A(�c	���W_U#�tr0���X���6���*4f'���������,�a�\�'��ؗ,�����������sP�w!���I��Ή������E������P��_W<t���j�tFt���򛤞��G�S�/>����ԝ�Έ~߈5RZ7%Gu�_�LKkÐ��4�{��E���,�﯅D���\<�xlܡm{�s}���!=��,-�n��`�.4�t���7u��P��OK싿�:��)؏��.	���8���	X�܇�7��t�箲��2�`0]Y΋�����:��	-�[���|тY?j��V#$8q/���O��^7�*��`�T�(�V��ŗN�Qt�;61���5���+�P3�Ns�9|iX,0w�3�����f7f"���G�^0fS֖?���͔u�duR�B�	�|���bc��W�I˂�,H�;�Ny��N�aKkO,�?a]�{� ^�N3���@����3�0^�Uptw�xsƄ��n���p܃��m��q�Y�����Ҝ�F-=�g'�Z��?c����]�@�7�䶬�vrk�^���'{����w��)�Ȝ��d�H��);�1���79-���^N��It7X�`g������yޘ�\���^��i�)�r��=y;rr�@���[xk�w�׉�JBMyD8��.�М��j`��Ԣ�Ʊ|W�Nc-�q\WFE�-�����)�W�b���Q?P��-zN�穲&�I���4�����2ԳBpD7]"�#�>����k҉�t���_sN.�����\�������uX�nQ��%�g�W9������C�W7�"K램NA8�?�N��uϝ�?��nЊ���x��H3:�[c�0�V��:@S`w�V�W�Z�!f�fV����Qvwb� $�sfŀ�w�o^2F�c��>�G�w��������Iޟ��{t�e�7������sW�>1�!$5�f�J��Z��F{Pd���/�<r(O�xp��u�U�ʄQ�{
 �m���^�=:�n?���J����)Z��b���e+���S��َ+(�D��w<��-��a�
�a���h|�>�e���B&��d�/F�:j��Ŵ������㲒?ܲQt����)��^B�9J@��W��!��֞��̐ �>ۈ�UŬ3u�$+A�1U+�	z!��Й��7s[��Z���wu\PZ�� �z�bV�걩�����rj�C"z\J�8/B�(����j�;$/�~��w�S���.�$��է��U��F��FC�"���2��h���� �,ln<FD!��\�ǭ�!K)j��\EL�J�G�cF���y�d�4��t0�q�8�0��4�"�F����g�ZIT���aM���E�x2��s�����Z��m`o���TsY9�	��j`����|�Ng��� Ճq�שZ���a��犁.���ҫk?.��|�N��mJ