��/  �K��7�o[q�"���~dcS$Sj|�s�n�^j�����h2Rgj���FQ
�F�GV����pxnwcA�H �E|�a���ww���d��{�~�ȝx�G��YŰ��vE��d2(��(>�E9�Q��%�b��IK��~��F cl86���nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n����D3ӡ���p"�pM�x �GIc�W�	� ��S�w��Jƙ�����O�A|$a�p(t�]7h����B�ړhb�Կ��v��Z�>կ䫒� ;�+�X���b������jTÿ*� r�f��T_�o����3	���O"��&����V�"%ΗD�����c��3��#|��B��
�,=$�%S^�EX:����v�P�.�s.��(�'�dF�A�4GgTu�j�"ed��GԞ3��:��C����К��n�*Y�6�kjz���J(O��_��`He�̟��	�"��zd��)�d�]�#�a���J������װ�\�p0U�ǈ5Xv i��Pr`�M�}�/�I
F͞R���ޛs:#xw�ܗY(��d~��Y�S�aW��.��+��O �ő��}T�֦��A#���Z�P��V�Ȗ!�w%Y���u*�e��c��~㐦 щb`W�r�#ov�4QŌox|���s�y�5Sp�1i��9�KGι����
�,�Ak"�#�Z��uO$/�r���u�U���ٔ�����A|[��Zͮ���\�a��b�Pf�E5��|�,5�6??�a"iTk�Â�]��+�|&p�[ #�����C����6�����a;�Ճ���ݎg���Ԓnz�o��+��Bb`N\��?�@J�ۗ
�̧��GZt���c�gX��Ym�Y#W�a,�H�tj�z�d̲c�Ȣ�Wvyk��w�x��+��K) �Le-Gl���r�6j�L˙�G%��a�/�*�ݻfz�^xt.M�����^�]CM�a'��c-1�o՗��hJ�����3��Nͻ��F�@�ܬ�T�(~8�S7��]J�2�MØN9�A �����F��z�T|p�q�)��@+��0]����Oz|��>?�u?��,gf����j'+N�/�!�����=��$mK!���6x}a�u뵺��/�w�_�����b�I�#ŧ,��*{�E�����O�f����7v���v9=�r��G^ai����`�JǱ�L@sQ�e�/� Xf��{btuPݖ��voZ&��9�d�[Ӆ9�űhE'R�ٲ�J�W��0�*�Ͱ�
��G"Ȋ��4�se]|� 2�v)+{�=Zr�/�1�ff�������j�����62�3䧛9V1�I�d_��d�w=�V�A
u��ؔ8��n�A/zz�%Y�?�-���z)k.m�ta{��D<e4�DK�b7<��sׁ��巻��8�(~*��U�����v^>JF�������t[gܽ>�l�
@ڷj�9UH�����1ri�f�w�s�)�O���7��z<j�A�W���Qr��pE:��L���?P��A���ѮB�t3� ��r�3+9������t��:�2�� SvJ���n���o!� 2�]}u�'��L���=1!��Ƞ�������͑�-���3��l������[v����h�م���)/��/r�7���nQT�NsP}F-!�]��
��[���%��A��^�z̀'o+)u5����^�"���4�w��ߏLęd;mm��G�y= D��ZM��ӷ���9�&HǃEG2`sKL6!p��*�V.ٔ�-v5[k��I9K�,�c�DRx,���X@#�"`Xs�ݿe!���]��J�R)VQ����Z�;����C��m#n�=kEX���rS����5/T�[#��4��e�5��K�:bӬ9�,5w��.��z����cC/Pk��)�E��M*iKC��o�.7U��S�{.���eU����*RS��Gb)*����j d��GWV��](�=)�{-7&lX���ݰ�z�0S��7U4�P�m��Xjs�	�e�kx��A9��6g�����1)6�L>48�b�]5f�Ȩ�Ϋ�ߺa˛Ur�^�V��$kVv7��l��R�����E
?�7s(m�=��R؆�p�.
,2�RpZ�:�1M���4ڨs�,tX/��?���у�kJD/�����~�*�F�Ư�[��|���)�o�V�n�xm�
����%���s��f�����F��=�jǟ�7��XǗ�7�R��o��=|o,ˮV�P�D)]��	D����6�p�����8a�)�dz��28RG�V��xÉT>%�y�>:�SŌ3��P� �;;�����b��Շ�y���q8B�#6�p������!�~��R��S�m��%��<���68mꞑc ��n�9X�v�t���<S�W�n.���D���5�$�y~��	:��}��_��>��G}�RxJ�@5j軷 S�Q9�̠l������wu�v����S�����i�7yc�����Q�����gz��hXp+��M�$�O���A�p�F�q�{�M�q�ք��?�+��9�p�Z����C�F�vqV=��!�\�o��.(.c��q�4����1�{+�6E'j2�ڣ���J�� �M����e�<�&h�˺vSCDE�����l�cDz�>~T�oy]�By1}kό�%��W2|:D7@Ѱ�o��l`�Eվ��z����OЎ���婮��0Cnw��#ø�j�0��"����\=�����:�=��$V��0P_�6��u����[ZbY���,��MW����ӒP�_�"��D<�L�V;��J�16
�i�����Ϩ��O�P����M	�7�HW�PЙ��d�*x	�! ���K~�b݈	�_���KHݏ#v����q�P $�M�	g=#��bm6cW��p�0�T��bu��?S�����=��¡�aE_2:�r6'�K[�#,�اJ�h9���'�Ȋ��J�m]o����eѲςy%��s����0�${l0��^t�v��'�����*%�tc�:���B"䊿CN�5�(֪��o�\g0&"s5��h5�a'U3DhWli���9��,�8�K� khn�z��#�%Q�6�Zx6��=��I������9V���mQ�n���5�λFd�_���W�g�����./���T�ɜl]�l��K!��� ���*<�D�zO�ƹ��hJ�J��y�I6���C��o<4m����f�o�+���v��������CI�\�
��>�9x�3==٤�8���$^�����n��#w��Y�G�<n	��H]p�"e�e"f����5��KL0J��^�o'#܎Y8�p=L<�D@m�$��X��=e���b��Mf��GW�T\����8(Ⱦ�/݀�}9�D��ez2s�)%3zez;�|%4���,�
	kq	�W���.Ї^�����|Rۏ�Z��r����&��ׁ�v��	��I�Z��>@�-��J~[�okq���4�+����!�Uׁ�k�PWʪt�Xm�� �FV>���6�*�F�;�/��۟�4�8�/�[aHXK�/���e��n���B�Y3�u��8[�a��J9��1�h���Ӹ��*�&8��!8�1��ב�R�h���cqj ����;�;��:Sv�3PŮ+p����&a��-�����bD^�߃�ߓ항��ˀC%2C����ΰ����ջ�K0`�aL��p�