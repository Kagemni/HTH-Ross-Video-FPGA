��/  =AA��j!&|�oo�N>��5/����K.\=��lV~��z0d�!�P���9�^}�*  ߌ<+����j[�z�_���o�h��g�X��[�	K��ִ�d�s��ƀy�d�������5�:���j�h�U.7I��p7�(G����I�����nhC_\��!ʝ��E}а9��z0�W@���W�&��}�PᵧIE�f�N��wX��u�ϛa�Ut10sAJ��ˌ%���n�n�W��ߌN��5=�8�:N|���gp�P�ظ��U��)�& g�J����[��kxO{F�D�P(X�i��q-�n��@ ۃE�ǚQ�(7��O�����g#��R�����KƤ��V�?�?�[��N���&L�,�0[D�*������iI�"<�� ���L0���I�R�d)�W�,5ǰ��t|
�.��x���#�۱��R�m�򓈛�d�����c�R��������k�/�~̀��#�q��.�~�8*#t�䊷ԊH�f+��i��,�r�x^/��m��$F�6�˪�6M�J$TH)44���|2�χ8 R y����H��uhe|/��u?�Z���\�*k�5m��Ίl��%Eq.������[r��=�0�����NC+ +1�lXK`�#%a>E�f���2�N��C�v=�MN��+p�b�Ǒ��L�f'�N*
:����{�A^���tu0QDJ�99��m��@"�c/ 	��l���l��@�2���l�\M���5�n����ص&�̐������
D;s��.��Dv�=�BY�+?���
hQ֯b%O�����l�:"��j���k��`"qުg`��ޝ�F���o���ܡ�n)�wwL,����JX�C�Nu�C�'r)��bz_Ųu�K���h: ���r\��P�iH ���.3��cDB�ڿ�<��CP����	<�g��O(����ض()(U�T�C����鑷��kr���T���Ӿ�[�޲�+�UN�3��gf5"���t����T_y<l�,���~/���C��?P˵N�HJ���de,&I~�d�z��=+�)��K̛18�q��4,1솦�C[< �>eY�;���Z+*Q���'�t'�h���A.��X@�g�{W����8��@↎C��\g�E��%8�f;���7�ڊ��j��c��bu�׎~B�<z�0�"&�k�Xu�&|L m���N.�ȢF�)fH�U�O�&P��Mie��,�?�o��`���pQ���6U��h�H���@0��`�]��PU�ahc�� �RF���iHǷ��Ȃ'���&�y(�����v-YPꦉQ�fE1V}���l[R��qԪ0��
�t�3R�x��%(B���O ��Ro���߹iD8��H�.�������> �h�t��}��Pn^�^M���řj5/I6�5�6:2�w�U�b(�B��CA�M(���ȆD��������$Hp�RR�I���~��Qpm��k�<?&01�X�����I�JKo�Oun�"�ǹ")�(%d^&m�U�e�X��i�O+�?��.y�9�'�YC!��5��9��ż�l粓���"d4��?|t��C�����nq_�L6�2�5�_�>���B�͖���܀�2A����%�SYt������sy���k�S��.���n΍#`oâ�Vͥ�L���Y��n�e�#Wzr��V9���p��8�>mׂ��r8�l9����0����8T�yY��CB��kX�6��[*���$�3����#���f5܄�M��p\'�E7�7���Ҵ��'2�`km��ѿ�Ӄ��l����u_�!+ua$�-�ʿ����8E���76��ЫȤUYE��R���O����k�K�L�$/�Y�w7V�y{ಇL�B�R�J��H�fMo��:��y�M&�^ѕ-���o�)���hP����y���%�������n5���E>Q+��~�:�+�&��"+`n���i"�
���ݨy�GHt�!�E��C���1,��&�&�!xטJ��^�)�� ��m��Բ��l��lDyOA��{�Y���P���U�4���.%ѽ��:\{��ʩ�P�E^$���U�|@*}�a%!�P�[�,���Sj����{�K-�|� ���0��v��H��xa͕�V������Z!~#*�{fw�~���ڕ�V��习g�����mt衇AJ�����]�-�� �:o_��f3��c����Ӆ�`��of��T5���w�K}�/���Z�c���Ίw&bH-^��T�����N�.�TA%ۥ+��D���u��+�fh�������2�s}�},+_�Ŏ�q�itT��SCW$�,͕,y/U��h�&\��{�r(S��RxЗtY\�!�		���FQC;��E'�Y{{y�]ݚ%����4���F&�� ��3Q�݅����u�1��L
}}�Kc~گ�Yc�hѠ�{c��v�>*�f��+�D�d+�)O�s!�;�&�,~���F��C�R����W�����	���\��_:ɹI��L��e2~�˂u���1���ǳ�R}�/�#�a��Q��;��7�,���@��J)<�e��,��C뇁�s�C���"��-�xl��ƺ]�J��H��D�G��y&�z[�f>k��?���`��/�P^7��a��u�I{�����������U��#`v��%^e��s�����p(�I��ߗ�v�;)�P��C��ꦡ"[